--Problem 5 TB
--All libraries in ModelSim default compile to work so we can access anything compiled under that library.
--No include managment, everything in the library you compile this to is automatically included.
--Use "compile to library" in ModelSim to pick where to compile
--I compiled all files to a folder called "Lab3" which is why I run
--library Lab3;
--use Problem5.all;