
module main(DATA_0_31,DATA_0_30,DATA_0_29,DATA_0_28,DATA_0_27,DATA_0_26,DATA_0_25,DATA_0_24,DATA_0_23,DATA_0_22,DATA_0_21,DATA_0_20,DATA_0_19,DATA_0_18,DATA_0_17,DATA_0_16,DATA_0_15,DATA_0_14,DATA_0_13,DATA_0_12,DATA_0_11,DATA_0_10,DATA_0_9,DATA_0_8,DATA_0_7,DATA_0_6,DATA_0_5,DATA_0_4,DATA_0_3,DATA_0_2,DATA_0_1,DATA_0_0,RESET,TM1,TM0,DATA_9_31,DATA_9_30,DATA_9_29,DATA_9_28,DATA_9_27,DATA_9_26,DATA_9_25,DATA_9_24,DATA_9_23,DATA_9_22,DATA_9_21,DATA_9_20,DATA_9_19,DATA_9_18,DATA_9_17,DATA_9_16,DATA_9_15,DATA_9_14,DATA_9_13,DATA_9_12,DATA_9_11,DATA_9_10,DATA_9_9,DATA_9_8,DATA_9_7,DATA_9_6,DATA_9_5,DATA_9_4,DATA_9_3,DATA_9_2,DATA_9_1,DATA_9_0,CRC_OUT_9_0,CRC_OUT_9_1,CRC_OUT_9_2,CRC_OUT_9_3,CRC_OUT_9_4,CRC_OUT_9_5,CRC_OUT_9_6,CRC_OUT_9_7,CRC_OUT_9_8,CRC_OUT_9_9,CRC_OUT_9_10,CRC_OUT_9_11,CRC_OUT_9_12,CRC_OUT_9_13,CRC_OUT_9_14,CRC_OUT_9_15,CRC_OUT_9_16,CRC_OUT_9_17,CRC_OUT_9_18,CRC_OUT_9_19,CRC_OUT_9_20,CRC_OUT_9_21,CRC_OUT_9_22,CRC_OUT_9_23,CRC_OUT_9_24,CRC_OUT_9_25,CRC_OUT_9_26,CRC_OUT_9_27,CRC_OUT_9_28,CRC_OUT_9_29,CRC_OUT_9_30,CRC_OUT_9_31,CRC_OUT_8_0,CRC_OUT_8_1,CRC_OUT_8_2,CRC_OUT_8_3,CRC_OUT_8_4,CRC_OUT_8_5,CRC_OUT_8_6,CRC_OUT_8_7,CRC_OUT_8_8,CRC_OUT_8_9,CRC_OUT_8_10,CRC_OUT_8_11,CRC_OUT_8_12,CRC_OUT_8_13,CRC_OUT_8_14,CRC_OUT_8_15,CRC_OUT_8_16,CRC_OUT_8_17,CRC_OUT_8_18,CRC_OUT_8_19,CRC_OUT_8_20,CRC_OUT_8_21,CRC_OUT_8_22,CRC_OUT_8_23,CRC_OUT_8_24,CRC_OUT_8_25,CRC_OUT_8_26,CRC_OUT_8_27,CRC_OUT_8_28,CRC_OUT_8_29,CRC_OUT_8_30,CRC_OUT_8_31,CRC_OUT_7_0,CRC_OUT_7_1,CRC_OUT_7_2,CRC_OUT_7_3,CRC_OUT_7_4,CRC_OUT_7_5,CRC_OUT_7_6,CRC_OUT_7_7,CRC_OUT_7_8,CRC_OUT_7_9,CRC_OUT_7_10,CRC_OUT_7_11,CRC_OUT_7_12,CRC_OUT_7_13,CRC_OUT_7_14,CRC_OUT_7_15,CRC_OUT_7_16,CRC_OUT_7_17,CRC_OUT_7_18,CRC_OUT_7_19,CRC_OUT_7_20,CRC_OUT_7_21,CRC_OUT_7_22,CRC_OUT_7_23,CRC_OUT_7_24,CRC_OUT_7_25,CRC_OUT_7_26,CRC_OUT_7_27,CRC_OUT_7_28,CRC_OUT_7_29,CRC_OUT_7_30,CRC_OUT_7_31,CRC_OUT_6_0,CRC_OUT_6_1,CRC_OUT_6_2,CRC_OUT_6_3,CRC_OUT_6_4,CRC_OUT_6_5,CRC_OUT_6_6,CRC_OUT_6_7,CRC_OUT_6_8,CRC_OUT_6_9,CRC_OUT_6_10,CRC_OUT_6_11,CRC_OUT_6_12,CRC_OUT_6_13,CRC_OUT_6_14,CRC_OUT_6_15,CRC_OUT_6_16,CRC_OUT_6_17,CRC_OUT_6_18,CRC_OUT_6_19,CRC_OUT_6_20,CRC_OUT_6_21,CRC_OUT_6_22,CRC_OUT_6_23,CRC_OUT_6_24,CRC_OUT_6_25,CRC_OUT_6_26,CRC_OUT_6_27,CRC_OUT_6_28,CRC_OUT_6_29,CRC_OUT_6_30,CRC_OUT_6_31,CRC_OUT_5_0,CRC_OUT_5_1,CRC_OUT_5_2,CRC_OUT_5_3,CRC_OUT_5_4,CRC_OUT_5_5,CRC_OUT_5_6,CRC_OUT_5_7,CRC_OUT_5_8,CRC_OUT_5_9,CRC_OUT_5_10,CRC_OUT_5_11,CRC_OUT_5_12,CRC_OUT_5_13,CRC_OUT_5_14,CRC_OUT_5_15,CRC_OUT_5_16,CRC_OUT_5_17,CRC_OUT_5_18,CRC_OUT_5_19,CRC_OUT_5_20,CRC_OUT_5_21,CRC_OUT_5_22,CRC_OUT_5_23,CRC_OUT_5_24,CRC_OUT_5_25,CRC_OUT_5_26,CRC_OUT_5_27,CRC_OUT_5_28,CRC_OUT_5_29,CRC_OUT_5_30,CRC_OUT_5_31,CRC_OUT_4_0,CRC_OUT_4_1,CRC_OUT_4_2,CRC_OUT_4_3,CRC_OUT_4_4,CRC_OUT_4_5,CRC_OUT_4_6,CRC_OUT_4_7,CRC_OUT_4_8,CRC_OUT_4_9,CRC_OUT_4_10,CRC_OUT_4_11,CRC_OUT_4_12,CRC_OUT_4_13,CRC_OUT_4_14,CRC_OUT_4_15,CRC_OUT_4_16,CRC_OUT_4_17,CRC_OUT_4_18,CRC_OUT_4_19,CRC_OUT_4_20,CRC_OUT_4_21,CRC_OUT_4_22,CRC_OUT_4_23,CRC_OUT_4_24,CRC_OUT_4_25,CRC_OUT_4_26,CRC_OUT_4_27,CRC_OUT_4_28,CRC_OUT_4_29,CRC_OUT_4_30,CRC_OUT_4_31,CRC_OUT_3_0,CRC_OUT_3_1,CRC_OUT_3_2,CRC_OUT_3_3,CRC_OUT_3_4,CRC_OUT_3_5,CRC_OUT_3_6,CRC_OUT_3_7,CRC_OUT_3_8,CRC_OUT_3_9,CRC_OUT_3_10,CRC_OUT_3_11,CRC_OUT_3_12,CRC_OUT_3_13,CRC_OUT_3_14,CRC_OUT_3_15,CRC_OUT_3_16,CRC_OUT_3_17,CRC_OUT_3_18,CRC_OUT_3_19,CRC_OUT_3_20,CRC_OUT_3_21,CRC_OUT_3_22,CRC_OUT_3_23,CRC_OUT_3_24,CRC_OUT_3_25,CRC_OUT_3_26,CRC_OUT_3_27,CRC_OUT_3_28,CRC_OUT_3_29,CRC_OUT_3_30,CRC_OUT_3_31,CRC_OUT_2_0,CRC_OUT_2_1,CRC_OUT_2_2,CRC_OUT_2_3,CRC_OUT_2_4,CRC_OUT_2_5,CRC_OUT_2_6,CRC_OUT_2_7,CRC_OUT_2_8,CRC_OUT_2_9,CRC_OUT_2_10,CRC_OUT_2_11,CRC_OUT_2_12,CRC_OUT_2_13,CRC_OUT_2_14,CRC_OUT_2_15,CRC_OUT_2_16,CRC_OUT_2_17,CRC_OUT_2_18,CRC_OUT_2_19,CRC_OUT_2_20,CRC_OUT_2_21,CRC_OUT_2_22,CRC_OUT_2_23,CRC_OUT_2_24,CRC_OUT_2_25,CRC_OUT_2_26,CRC_OUT_2_27,CRC_OUT_2_28,CRC_OUT_2_29,CRC_OUT_2_30,CRC_OUT_2_31,CRC_OUT_1_0,CRC_OUT_1_1,CRC_OUT_1_2,CRC_OUT_1_3,CRC_OUT_1_4,CRC_OUT_1_5,CRC_OUT_1_6,CRC_OUT_1_7,CRC_OUT_1_8,CRC_OUT_1_9,CRC_OUT_1_10,CRC_OUT_1_11,CRC_OUT_1_12,CRC_OUT_1_13,CRC_OUT_1_14,CRC_OUT_1_15,CRC_OUT_1_16,CRC_OUT_1_17,CRC_OUT_1_18,CRC_OUT_1_19,CRC_OUT_1_20,CRC_OUT_1_21,CRC_OUT_1_22,CRC_OUT_1_23,CRC_OUT_1_24,CRC_OUT_1_25,CRC_OUT_1_26,CRC_OUT_1_27,CRC_OUT_1_28,CRC_OUT_1_29,CRC_OUT_1_30,CRC_OUT_1_31);

input DATA_0_31;
input DATA_0_30;
input DATA_0_29;
input DATA_0_28;
input DATA_0_27;
input DATA_0_26;
input DATA_0_25;
input DATA_0_24;
input DATA_0_23;
input DATA_0_22;
input DATA_0_21;
input DATA_0_20;
input DATA_0_19;
input DATA_0_18;
input DATA_0_17;
input DATA_0_16;
input DATA_0_15;
input DATA_0_14;
input DATA_0_13;
input DATA_0_12;
input DATA_0_11;
input DATA_0_10;
input DATA_0_9;
input DATA_0_8;
input DATA_0_7;
input DATA_0_6;
input DATA_0_5;
input DATA_0_4;
input DATA_0_3;
input DATA_0_2;
input DATA_0_1;
input DATA_0_0;
input RESET;
input TM1;
input TM0;

output DATA_9_31;
output DATA_9_30;
output DATA_9_29;
output DATA_9_28;
output DATA_9_27;
output DATA_9_26;
output DATA_9_25;
output DATA_9_24;
output DATA_9_23;
output DATA_9_22;
output DATA_9_21;
output DATA_9_20;
output DATA_9_19;
output DATA_9_18;
output DATA_9_17;
output DATA_9_16;
output DATA_9_15;
output DATA_9_14;
output DATA_9_13;
output DATA_9_12;
output DATA_9_11;
output DATA_9_10;
output DATA_9_9;
output DATA_9_8;
output DATA_9_7;
output DATA_9_6;
output DATA_9_5;
output DATA_9_4;
output DATA_9_3;
output DATA_9_2;
output DATA_9_1;
output DATA_9_0;
output CRC_OUT_9_0;
output CRC_OUT_9_1;
output CRC_OUT_9_2;
output CRC_OUT_9_3;
output CRC_OUT_9_4;
output CRC_OUT_9_5;
output CRC_OUT_9_6;
output CRC_OUT_9_7;
output CRC_OUT_9_8;
output CRC_OUT_9_9;
output CRC_OUT_9_10;
output CRC_OUT_9_11;
output CRC_OUT_9_12;
output CRC_OUT_9_13;
output CRC_OUT_9_14;
output CRC_OUT_9_15;
output CRC_OUT_9_16;
output CRC_OUT_9_17;
output CRC_OUT_9_18;
output CRC_OUT_9_19;
output CRC_OUT_9_20;
output CRC_OUT_9_21;
output CRC_OUT_9_22;
output CRC_OUT_9_23;
output CRC_OUT_9_24;
output CRC_OUT_9_25;
output CRC_OUT_9_26;
output CRC_OUT_9_27;
output CRC_OUT_9_28;
output CRC_OUT_9_29;
output CRC_OUT_9_30;
output CRC_OUT_9_31;
output CRC_OUT_8_0;
output CRC_OUT_8_1;
output CRC_OUT_8_2;
output CRC_OUT_8_3;
output CRC_OUT_8_4;
output CRC_OUT_8_5;
output CRC_OUT_8_6;
output CRC_OUT_8_7;
output CRC_OUT_8_8;
output CRC_OUT_8_9;
output CRC_OUT_8_10;
output CRC_OUT_8_11;
output CRC_OUT_8_12;
output CRC_OUT_8_13;
output CRC_OUT_8_14;
output CRC_OUT_8_15;
output CRC_OUT_8_16;
output CRC_OUT_8_17;
output CRC_OUT_8_18;
output CRC_OUT_8_19;
output CRC_OUT_8_20;
output CRC_OUT_8_21;
output CRC_OUT_8_22;
output CRC_OUT_8_23;
output CRC_OUT_8_24;
output CRC_OUT_8_25;
output CRC_OUT_8_26;
output CRC_OUT_8_27;
output CRC_OUT_8_28;
output CRC_OUT_8_29;
output CRC_OUT_8_30;
output CRC_OUT_8_31;
output CRC_OUT_7_0;
output CRC_OUT_7_1;
output CRC_OUT_7_2;
output CRC_OUT_7_3;
output CRC_OUT_7_4;
output CRC_OUT_7_5;
output CRC_OUT_7_6;
output CRC_OUT_7_7;
output CRC_OUT_7_8;
output CRC_OUT_7_9;
output CRC_OUT_7_10;
output CRC_OUT_7_11;
output CRC_OUT_7_12;
output CRC_OUT_7_13;
output CRC_OUT_7_14;
output CRC_OUT_7_15;
output CRC_OUT_7_16;
output CRC_OUT_7_17;
output CRC_OUT_7_18;
output CRC_OUT_7_19;
output CRC_OUT_7_20;
output CRC_OUT_7_21;
output CRC_OUT_7_22;
output CRC_OUT_7_23;
output CRC_OUT_7_24;
output CRC_OUT_7_25;
output CRC_OUT_7_26;
output CRC_OUT_7_27;
output CRC_OUT_7_28;
output CRC_OUT_7_29;
output CRC_OUT_7_30;
output CRC_OUT_7_31;
output CRC_OUT_6_0;
output CRC_OUT_6_1;
output CRC_OUT_6_2;
output CRC_OUT_6_3;
output CRC_OUT_6_4;
output CRC_OUT_6_5;
output CRC_OUT_6_6;
output CRC_OUT_6_7;
output CRC_OUT_6_8;
output CRC_OUT_6_9;
output CRC_OUT_6_10;
output CRC_OUT_6_11;
output CRC_OUT_6_12;
output CRC_OUT_6_13;
output CRC_OUT_6_14;
output CRC_OUT_6_15;
output CRC_OUT_6_16;
output CRC_OUT_6_17;
output CRC_OUT_6_18;
output CRC_OUT_6_19;
output CRC_OUT_6_20;
output CRC_OUT_6_21;
output CRC_OUT_6_22;
output CRC_OUT_6_23;
output CRC_OUT_6_24;
output CRC_OUT_6_25;
output CRC_OUT_6_26;
output CRC_OUT_6_27;
output CRC_OUT_6_28;
output CRC_OUT_6_29;
output CRC_OUT_6_30;
output CRC_OUT_6_31;
output CRC_OUT_5_0;
output CRC_OUT_5_1;
output CRC_OUT_5_2;
output CRC_OUT_5_3;
output CRC_OUT_5_4;
output CRC_OUT_5_5;
output CRC_OUT_5_6;
output CRC_OUT_5_7;
output CRC_OUT_5_8;
output CRC_OUT_5_9;
output CRC_OUT_5_10;
output CRC_OUT_5_11;
output CRC_OUT_5_12;
output CRC_OUT_5_13;
output CRC_OUT_5_14;
output CRC_OUT_5_15;
output CRC_OUT_5_16;
output CRC_OUT_5_17;
output CRC_OUT_5_18;
output CRC_OUT_5_19;
output CRC_OUT_5_20;
output CRC_OUT_5_21;
output CRC_OUT_5_22;
output CRC_OUT_5_23;
output CRC_OUT_5_24;
output CRC_OUT_5_25;
output CRC_OUT_5_26;
output CRC_OUT_5_27;
output CRC_OUT_5_28;
output CRC_OUT_5_29;
output CRC_OUT_5_30;
output CRC_OUT_5_31;
output CRC_OUT_4_0;
output CRC_OUT_4_1;
output CRC_OUT_4_2;
output CRC_OUT_4_3;
output CRC_OUT_4_4;
output CRC_OUT_4_5;
output CRC_OUT_4_6;
output CRC_OUT_4_7;
output CRC_OUT_4_8;
output CRC_OUT_4_9;
output CRC_OUT_4_10;
output CRC_OUT_4_11;
output CRC_OUT_4_12;
output CRC_OUT_4_13;
output CRC_OUT_4_14;
output CRC_OUT_4_15;
output CRC_OUT_4_16;
output CRC_OUT_4_17;
output CRC_OUT_4_18;
output CRC_OUT_4_19;
output CRC_OUT_4_20;
output CRC_OUT_4_21;
output CRC_OUT_4_22;
output CRC_OUT_4_23;
output CRC_OUT_4_24;
output CRC_OUT_4_25;
output CRC_OUT_4_26;
output CRC_OUT_4_27;
output CRC_OUT_4_28;
output CRC_OUT_4_29;
output CRC_OUT_4_30;
output CRC_OUT_4_31;
output CRC_OUT_3_0;
output CRC_OUT_3_1;
output CRC_OUT_3_2;
output CRC_OUT_3_3;
output CRC_OUT_3_4;
output CRC_OUT_3_5;
output CRC_OUT_3_6;
output CRC_OUT_3_7;
output CRC_OUT_3_8;
output CRC_OUT_3_9;
output CRC_OUT_3_10;
output CRC_OUT_3_11;
output CRC_OUT_3_12;
output CRC_OUT_3_13;
output CRC_OUT_3_14;
output CRC_OUT_3_15;
output CRC_OUT_3_16;
output CRC_OUT_3_17;
output CRC_OUT_3_18;
output CRC_OUT_3_19;
output CRC_OUT_3_20;
output CRC_OUT_3_21;
output CRC_OUT_3_22;
output CRC_OUT_3_23;
output CRC_OUT_3_24;
output CRC_OUT_3_25;
output CRC_OUT_3_26;
output CRC_OUT_3_27;
output CRC_OUT_3_28;
output CRC_OUT_3_29;
output CRC_OUT_3_30;
output CRC_OUT_3_31;
output CRC_OUT_2_0;
output CRC_OUT_2_1;
output CRC_OUT_2_2;
output CRC_OUT_2_3;
output CRC_OUT_2_4;
output CRC_OUT_2_5;
output CRC_OUT_2_6;
output CRC_OUT_2_7;
output CRC_OUT_2_8;
output CRC_OUT_2_9;
output CRC_OUT_2_10;
output CRC_OUT_2_11;
output CRC_OUT_2_12;
output CRC_OUT_2_13;
output CRC_OUT_2_14;
output CRC_OUT_2_15;
output CRC_OUT_2_16;
output CRC_OUT_2_17;
output CRC_OUT_2_18;
output CRC_OUT_2_19;
output CRC_OUT_2_20;
output CRC_OUT_2_21;
output CRC_OUT_2_22;
output CRC_OUT_2_23;
output CRC_OUT_2_24;
output CRC_OUT_2_25;
output CRC_OUT_2_26;
output CRC_OUT_2_27;
output CRC_OUT_2_28;
output CRC_OUT_2_29;
output CRC_OUT_2_30;
output CRC_OUT_2_31;
output CRC_OUT_1_0;
output CRC_OUT_1_1;
output CRC_OUT_1_2;
output CRC_OUT_1_3;
output CRC_OUT_1_4;
output CRC_OUT_1_5;
output CRC_OUT_1_6;
output CRC_OUT_1_7;
output CRC_OUT_1_8;
output CRC_OUT_1_9;
output CRC_OUT_1_10;
output CRC_OUT_1_11;
output CRC_OUT_1_12;
output CRC_OUT_1_13;
output CRC_OUT_1_14;
output CRC_OUT_1_15;
output CRC_OUT_1_16;
output CRC_OUT_1_17;
output CRC_OUT_1_18;
output CRC_OUT_1_19;
output CRC_OUT_1_20;
output CRC_OUT_1_21;
output CRC_OUT_1_22;
output CRC_OUT_1_23;
output CRC_OUT_1_24;
output CRC_OUT_1_25;
output CRC_OUT_1_26;
output CRC_OUT_1_27;
output CRC_OUT_1_28;
output CRC_OUT_1_29;
output CRC_OUT_1_30;
output CRC_OUT_1_31;
//There are problems because CRC out is declared as an output and a wire.
wire 	WX485,WX487,WX489,WX491,WX493,WX495,WX497
	,WX499,WX501,WX503,WX505,WX507,WX509,WX511,WX513
	,WX515,WX517,WX519,WX521,WX523,WX525,WX527,WX529
	,WX531,WX533,WX535,WX537,WX539,WX541,WX543,WX545
	,WX547,WX645,WX647,WX649,WX651,WX653,WX655,WX657
	,WX659,WX661,WX663,WX665,WX667,WX669,WX671,WX673
	,WX675,WX677,WX679,WX681,WX683,WX685,WX687,WX689
	,WX691,WX693,WX695,WX697,WX699,WX701,WX703,WX705
	,WX707,WX709,WX711,WX713,WX715,WX717,WX719,WX721
	,WX723,WX725,WX727,WX729,WX731,WX733,WX735,WX737
	,WX739,WX741,WX743,WX745,WX747,WX749,WX751,WX753
	,WX755,WX757,WX759,WX761,WX763,WX765,WX767,WX769
	,WX771,WX773,WX775,WX777,WX779,WX781,WX783,WX785
	,WX787,WX789,WX791,WX793,WX795,WX797,WX799,WX801
	,WX803,WX805,WX807,WX809,WX811,WX813,WX815,WX817
	,WX819,WX821,WX823,WX825,WX827,WX829,WX831,WX833
	,WX835,WX837,WX839,WX841,WX843,WX845,WX847,WX849
	,WX851,WX853,WX855,WX857,WX859,WX861,WX863,WX865
	,WX867,WX869,WX871,WX873,WX875,WX877,WX879,WX881
	,WX883,WX885,WX887,WX889,WX891,WX893,WX895,WX897
	,WX899,WX1778,WX1780,WX1782,WX1784,WX1786,WX1788,WX1790
	,WX1792,WX1794,WX1796,WX1798,WX1800,WX1802,WX1804,WX1806
	,WX1808,WX1810,WX1812,WX1814,WX1816,WX1818,WX1820,WX1822
	,WX1824,WX1826,WX1828,WX1830,WX1832,WX1834,WX1836,WX1838
	,WX1840,WX1938,WX1940,WX1942,WX1944,WX1946,WX1948,WX1950
	,WX1952,WX1954,WX1956,WX1958,WX1960,WX1962,WX1964,WX1966
	,WX1968,WX1970,WX1972,WX1974,WX1976,WX1978,WX1980,WX1982
	,WX1984,WX1986,WX1988,WX1990,WX1992,WX1994,WX1996,WX1998
	,WX2000,WX2002,WX2004,WX2006,WX2008,WX2010,WX2012,WX2014
	,WX2016,WX2018,WX2020,WX2022,WX2024,WX2026,WX2028,WX2030
	,WX2032,WX2034,WX2036,WX2038,WX2040,WX2042,WX2044,WX2046
	,WX2048,WX2050,WX2052,WX2054,WX2056,WX2058,WX2060,WX2062
	,WX2064,WX2066,WX2068,WX2070,WX2072,WX2074,WX2076,WX2078
	,WX2080,WX2082,WX2084,WX2086,WX2088,WX2090,WX2092,WX2094
	,WX2096,WX2098,WX2100,WX2102,WX2104,WX2106,WX2108,WX2110
	,WX2112,WX2114,WX2116,WX2118,WX2120,WX2122,WX2124,WX2126
	,WX2128,WX2130,WX2132,WX2134,WX2136,WX2138,WX2140,WX2142
	,WX2144,WX2146,WX2148,WX2150,WX2152,WX2154,WX2156,WX2158
	,WX2160,WX2162,WX2164,WX2166,WX2168,WX2170,WX2172,WX2174
	,WX2176,WX2178,WX2180,WX2182,WX2184,WX2186,WX2188,WX2190
	,WX2192,WX3071,WX3073,WX3075,WX3077,WX3079,WX3081,WX3083
	,WX3085,WX3087,WX3089,WX3091,WX3093,WX3095,WX3097,WX3099
	,WX3101,WX3103,WX3105,WX3107,WX3109,WX3111,WX3113,WX3115
	,WX3117,WX3119,WX3121,WX3123,WX3125,WX3127,WX3129,WX3131
	,WX3133,WX3231,WX3233,WX3235,WX3237,WX3239,WX3241,WX3243
	,WX3245,WX3247,WX3249,WX3251,WX3253,WX3255,WX3257,WX3259
	,WX3261,WX3263,WX3265,WX3267,WX3269,WX3271,WX3273,WX3275
	,WX3277,WX3279,WX3281,WX3283,WX3285,WX3287,WX3289,WX3291
	,WX3293,WX3295,WX3297,WX3299,WX3301,WX3303,WX3305,WX3307
	,WX3309,WX3311,WX3313,WX3315,WX3317,WX3319,WX3321,WX3323
	,WX3325,WX3327,WX3329,WX3331,WX3333,WX3335,WX3337,WX3339
	,WX3341,WX3343,WX3345,WX3347,WX3349,WX3351,WX3353,WX3355
	,WX3357,WX3359,WX3361,WX3363,WX3365,WX3367,WX3369,WX3371
	,WX3373,WX3375,WX3377,WX3379,WX3381,WX3383,WX3385,WX3387
	,WX3389,WX3391,WX3393,WX3395,WX3397,WX3399,WX3401,WX3403
	,WX3405,WX3407,WX3409,WX3411,WX3413,WX3415,WX3417,WX3419
	,WX3421,WX3423,WX3425,WX3427,WX3429,WX3431,WX3433,WX3435
	,WX3437,WX3439,WX3441,WX3443,WX3445,WX3447,WX3449,WX3451
	,WX3453,WX3455,WX3457,WX3459,WX3461,WX3463,WX3465,WX3467
	,WX3469,WX3471,WX3473,WX3475,WX3477,WX3479,WX3481,WX3483
	,WX3485,WX4364,WX4366,WX4368,WX4370,WX4372,WX4374,WX4376
	,WX4378,WX4380,WX4382,WX4384,WX4386,WX4388,WX4390,WX4392
	,WX4394,WX4396,WX4398,WX4400,WX4402,WX4404,WX4406,WX4408
	,WX4410,WX4412,WX4414,WX4416,WX4418,WX4420,WX4422,WX4424
	,WX4426,WX4524,WX4526,WX4528,WX4530,WX4532,WX4534,WX4536
	,WX4538,WX4540,WX4542,WX4544,WX4546,WX4548,WX4550,WX4552
	,WX4554,WX4556,WX4558,WX4560,WX4562,WX4564,WX4566,WX4568
	,WX4570,WX4572,WX4574,WX4576,WX4578,WX4580,WX4582,WX4584
	,WX4586,WX4588,WX4590,WX4592,WX4594,WX4596,WX4598,WX4600
	,WX4602,WX4604,WX4606,WX4608,WX4610,WX4612,WX4614,WX4616
	,WX4618,WX4620,WX4622,WX4624,WX4626,WX4628,WX4630,WX4632
	,WX4634,WX4636,WX4638,WX4640,WX4642,WX4644,WX4646,WX4648
	,WX4650,WX4652,WX4654,WX4656,WX4658,WX4660,WX4662,WX4664
	,WX4666,WX4668,WX4670,WX4672,WX4674,WX4676,WX4678,WX4680
	,WX4682,WX4684,WX4686,WX4688,WX4690,WX4692,WX4694,WX4696
	,WX4698,WX4700,WX4702,WX4704,WX4706,WX4708,WX4710,WX4712
	,WX4714,WX4716,WX4718,WX4720,WX4722,WX4724,WX4726,WX4728
	,WX4730,WX4732,WX4734,WX4736,WX4738,WX4740,WX4742,WX4744
	,WX4746,WX4748,WX4750,WX4752,WX4754,WX4756,WX4758,WX4760
	,WX4762,WX4764,WX4766,WX4768,WX4770,WX4772,WX4774,WX4776
	,WX4778,WX5657,WX5659,WX5661,WX5663,WX5665,WX5667,WX5669
	,WX5671,WX5673,WX5675,WX5677,WX5679,WX5681,WX5683,WX5685
	,WX5687,WX5689,WX5691,WX5693,WX5695,WX5697,WX5699,WX5701
	,WX5703,WX5705,WX5707,WX5709,WX5711,WX5713,WX5715,WX5717
	,WX5719,WX5817,WX5819,WX5821,WX5823,WX5825,WX5827,WX5829
	,WX5831,WX5833,WX5835,WX5837,WX5839,WX5841,WX5843,WX5845
	,WX5847,WX5849,WX5851,WX5853,WX5855,WX5857,WX5859,WX5861
	,WX5863,WX5865,WX5867,WX5869,WX5871,WX5873,WX5875,WX5877
	,WX5879,WX5881,WX5883,WX5885,WX5887,WX5889,WX5891,WX5893
	,WX5895,WX5897,WX5899,WX5901,WX5903,WX5905,WX5907,WX5909
	,WX5911,WX5913,WX5915,WX5917,WX5919,WX5921,WX5923,WX5925
	,WX5927,WX5929,WX5931,WX5933,WX5935,WX5937,WX5939,WX5941
	,WX5943,WX5945,WX5947,WX5949,WX5951,WX5953,WX5955,WX5957
	,WX5959,WX5961,WX5963,WX5965,WX5967,WX5969,WX5971,WX5973
	,WX5975,WX5977,WX5979,WX5981,WX5983,WX5985,WX5987,WX5989
	,WX5991,WX5993,WX5995,WX5997,WX5999,WX6001,WX6003,WX6005
	,WX6007,WX6009,WX6011,WX6013,WX6015,WX6017,WX6019,WX6021
	,WX6023,WX6025,WX6027,WX6029,WX6031,WX6033,WX6035,WX6037
	,WX6039,WX6041,WX6043,WX6045,WX6047,WX6049,WX6051,WX6053
	,WX6055,WX6057,WX6059,WX6061,WX6063,WX6065,WX6067,WX6069
	,WX6071,WX6950,WX6952,WX6954,WX6956,WX6958,WX6960,WX6962
	,WX6964,WX6966,WX6968,WX6970,WX6972,WX6974,WX6976,WX6978
	,WX6980,WX6982,WX6984,WX6986,WX6988,WX6990,WX6992,WX6994
	,WX6996,WX6998,WX7000,WX7002,WX7004,WX7006,WX7008,WX7010
	,WX7012,WX7110,WX7112,WX7114,WX7116,WX7118,WX7120,WX7122
	,WX7124,WX7126,WX7128,WX7130,WX7132,WX7134,WX7136,WX7138
	,WX7140,WX7142,WX7144,WX7146,WX7148,WX7150,WX7152,WX7154
	,WX7156,WX7158,WX7160,WX7162,WX7164,WX7166,WX7168,WX7170
	,WX7172,WX7174,WX7176,WX7178,WX7180,WX7182,WX7184,WX7186
	,WX7188,WX7190,WX7192,WX7194,WX7196,WX7198,WX7200,WX7202
	,WX7204,WX7206,WX7208,WX7210,WX7212,WX7214,WX7216,WX7218
	,WX7220,WX7222,WX7224,WX7226,WX7228,WX7230,WX7232,WX7234
	,WX7236,WX7238,WX7240,WX7242,WX7244,WX7246,WX7248,WX7250
	,WX7252,WX7254,WX7256,WX7258,WX7260,WX7262,WX7264,WX7266
	,WX7268,WX7270,WX7272,WX7274,WX7276,WX7278,WX7280,WX7282
	,WX7284,WX7286,WX7288,WX7290,WX7292,WX7294,WX7296,WX7298
	,WX7300,WX7302,WX7304,WX7306,WX7308,WX7310,WX7312,WX7314
	,WX7316,WX7318,WX7320,WX7322,WX7324,WX7326,WX7328,WX7330
	,WX7332,WX7334,WX7336,WX7338,WX7340,WX7342,WX7344,WX7346
	,WX7348,WX7350,WX7352,WX7354,WX7356,WX7358,WX7360,WX7362
	,WX7364,WX8243,WX8245,WX8247,WX8249,WX8251,WX8253,WX8255
	,WX8257,WX8259,WX8261,WX8263,WX8265,WX8267,WX8269,WX8271
	,WX8273,WX8275,WX8277,WX8279,WX8281,WX8283,WX8285,WX8287
	,WX8289,WX8291,WX8293,WX8295,WX8297,WX8299,WX8301,WX8303
	,WX8305,WX8403,WX8405,WX8407,WX8409,WX8411,WX8413,WX8415
	,WX8417,WX8419,WX8421,WX8423,WX8425,WX8427,WX8429,WX8431
	,WX8433,WX8435,WX8437,WX8439,WX8441,WX8443,WX8445,WX8447
	,WX8449,WX8451,WX8453,WX8455,WX8457,WX8459,WX8461,WX8463
	,WX8465,WX8467,WX8469,WX8471,WX8473,WX8475,WX8477,WX8479
	,WX8481,WX8483,WX8485,WX8487,WX8489,WX8491,WX8493,WX8495
	,WX8497,WX8499,WX8501,WX8503,WX8505,WX8507,WX8509,WX8511
	,WX8513,WX8515,WX8517,WX8519,WX8521,WX8523,WX8525,WX8527
	,WX8529,WX8531,WX8533,WX8535,WX8537,WX8539,WX8541,WX8543
	,WX8545,WX8547,WX8549,WX8551,WX8553,WX8555,WX8557,WX8559
	,WX8561,WX8563,WX8565,WX8567,WX8569,WX8571,WX8573,WX8575
	,WX8577,WX8579,WX8581,WX8583,WX8585,WX8587,WX8589,WX8591
	,WX8593,WX8595,WX8597,WX8599,WX8601,WX8603,WX8605,WX8607
	,WX8609,WX8611,WX8613,WX8615,WX8617,WX8619,WX8621,WX8623
	,WX8625,WX8627,WX8629,WX8631,WX8633,WX8635,WX8637,WX8639
	,WX8641,WX8643,WX8645,WX8647,WX8649,WX8651,WX8653,WX8655
	,WX8657,WX9536,WX9538,WX9540,WX9542,WX9544,WX9546,WX9548
	,WX9550,WX9552,WX9554,WX9556,WX9558,WX9560,WX9562,WX9564
	,WX9566,WX9568,WX9570,WX9572,WX9574,WX9576,WX9578,WX9580
	,WX9582,WX9584,WX9586,WX9588,WX9590,WX9592,WX9594,WX9596
	,WX9598,WX9696,WX9698,WX9700,WX9702,WX9704,WX9706,WX9708
	,WX9710,WX9712,WX9714,WX9716,WX9718,WX9720,WX9722,WX9724
	,WX9726,WX9728,WX9730,WX9732,WX9734,WX9736,WX9738,WX9740
	,WX9742,WX9744,WX9746,WX9748,WX9750,WX9752,WX9754,WX9756
	,WX9758,WX9760,WX9762,WX9764,WX9766,WX9768,WX9770,WX9772
	,WX9774,WX9776,WX9778,WX9780,WX9782,WX9784,WX9786,WX9788
	,WX9790,WX9792,WX9794,WX9796,WX9798,WX9800,WX9802,WX9804
	,WX9806,WX9808,WX9810,WX9812,WX9814,WX9816,WX9818,WX9820
	,WX9822,WX9824,WX9826,WX9828,WX9830,WX9832,WX9834,WX9836
	,WX9838,WX9840,WX9842,WX9844,WX9846,WX9848,WX9850,WX9852
	,WX9854,WX9856,WX9858,WX9860,WX9862,WX9864,WX9866,WX9868
	,WX9870,WX9872,WX9874,WX9876,WX9878,WX9880,WX9882,WX9884
	,WX9886,WX9888,WX9890,WX9892,WX9894,WX9896,WX9898,WX9900
	,WX9902,WX9904,WX9906,WX9908,WX9910,WX9912,WX9914,WX9916
	,WX9918,WX9920,WX9922,WX9924,WX9926,WX9928,WX9930,WX9932
	,WX9934,WX9936,WX9938,WX9940,WX9942,WX9944,WX9946,WX9948
	,WX9950,WX10829,WX10831,WX10833,WX10835,WX10837,WX10839,WX10841
	,WX10843,WX10845,WX10847,WX10849,WX10851,WX10853,WX10855,WX10857
	,WX10859,WX10861,WX10863,WX10865,WX10867,WX10869,WX10871,WX10873
	,WX10875,WX10877,WX10879,WX10881,WX10883,WX10885,WX10887,WX10889
	,WX10891,WX10989,WX10991,WX10993,WX10995,WX10997,WX10999,WX11001
	,WX11003,WX11005,WX11007,WX11009,WX11011,WX11013,WX11015,WX11017
	,WX11019,WX11021,WX11023,WX11025,WX11027,WX11029,WX11031,WX11033
	,WX11035,WX11037,WX11039,WX11041,WX11043,WX11045,WX11047,WX11049
	,WX11051,WX11053,WX11055,WX11057,WX11059,WX11061,WX11063,WX11065
	,WX11067,WX11069,WX11071,WX11073,WX11075,WX11077,WX11079,WX11081
	,WX11083,WX11085,WX11087,WX11089,WX11091,WX11093,WX11095,WX11097
	,WX11099,WX11101,WX11103,WX11105,WX11107,WX11109,WX11111,WX11113
	,WX11115,WX11117,WX11119,WX11121,WX11123,WX11125,WX11127,WX11129
	,WX11131,WX11133,WX11135,WX11137,WX11139,WX11141,WX11143,WX11145
	,WX11147,WX11149,WX11151,WX11153,WX11155,WX11157,WX11159,WX11161
	,WX11163,WX11165,WX11167,WX11169,WX11171,WX11173,WX11175,WX11177
	,WX11179,WX11181,WX11183,WX11185,WX11187,WX11189,WX11191,WX11193
	,WX11195,WX11197,WX11199,WX11201,WX11203,WX11205,WX11207,WX11209
	,WX11211,WX11213,WX11215,WX11217,WX11219,WX11221,WX11223,WX11225
	,WX11227,WX11229,WX11231,WX11233,WX11235,WX11237,WX11239,WX11241
	,WX11243,WX11574,WX10281,WX8988,WX7695,WX6402,WX5109,WX3816
	,WX2523,WX1230,WX11344,WX11343,WX10051,WX10050,WX8758,WX8757
	,WX7465,WX7464,WX6172,WX6171,WX4879,WX4878,WX3586,WX3585
	,WX2293,WX2292,WX1000,WX999,WX11342,WX11341,WX11340,WX10049
	,WX10048,WX10047,WX8756,WX8755,WX8754,WX7463,WX7462,WX7461
	,WX6170,WX6169,WX6168,WX4877,WX4876,WX4875,WX3584,WX3583
	,WX3582,WX2291,WX2290,WX2289,WX998,WX997,WX996,WX1005
	,WX1004,WX1002,WX2298,WX2297,WX2295,WX3591,WX3590,WX3588
	,WX4884,WX4883,WX4881,WX6177,WX6176,WX6174,WX7470,WX7469
	,WX7467,WX8763,WX8762,WX8760,WX10056,WX10055,WX10053,WX11349
	,WX11348,WX11346,WX1003,WX1001,WX2296,WX2294,WX3589,WX3587
	,WX4882,WX4880,WX6175,WX6173,WX7468,WX7466,WX8761,WX8759
	,WX10054,WX10052,WX11347,WX11345,WX1263,WX2556,WX3849,WX5142
	,WX6435,WX7728,WX9021,WX10314,WX11607,WX11242,WX11240,WX11238
	,WX11236,WX11234,WX11232,WX11230,WX11228,WX11226,WX11224,WX11222
	,WX11220,WX11218,WX11216,WX11214,WX11212,WX11210,WX11208,WX11206
	,WX11204,WX11202,WX11200,WX11198,WX11196,WX11194,WX11192,WX11190
	,WX11188,WX11186,WX11184,WX11182,WX11180,WX11178,WX11176,WX11174
	,WX11172,WX11170,WX11168,WX11166,WX11164,WX11162,WX11160,WX11158
	,WX11156,WX11154,WX11152,WX11150,WX11148,WX11146,WX11144,WX11142
	,WX11140,WX11138,WX11136,WX11134,WX11132,WX11130,WX11128,WX11126
	,WX11124,WX11122,WX11120,WX11118,WX11116,WX11114,WX11112,WX11110
	,WX11108,WX11106,WX11104,WX11102,WX11100,WX11098,WX11096,WX11094
	,WX11092,WX11090,WX11088,WX11086,WX11084,WX11082,WX11080,WX11078
	,WX11076,WX11074,WX11072,WX11070,WX11068,WX11066,WX11064,WX11062
	,WX11060,WX11058,WX11056,WX11054,WX11052,WX10888,WX10886,WX10884
	,WX10882,WX10880,WX10878,WX10876,WX10874,WX10872,WX10870,WX10868
	,WX10866,WX10864,WX10862,WX10860,WX10858,WX10856,WX10854,WX10852
	,WX10850,WX10848,WX10846,WX10844,WX10842,WX10840,WX10838,WX10836
	,WX10834,WX10832,WX10830,WX10828,WX9949,WX9947,WX9945,WX9943
	,WX9941,WX9939,WX9937,WX9935,WX9933,WX9931,WX9929,WX9927
	,WX9925,WX9923,WX9921,WX9919,WX9917,WX9915,WX9913,WX9911
	,WX9909,WX9907,WX9905,WX9903,WX9901,WX9899,WX9897,WX9895
	,WX9893,WX9891,WX9889,WX9887,WX9885,WX9883,WX9881,WX9879
	,WX9877,WX9875,WX9873,WX9871,WX9869,WX9867,WX9865,WX9863
	,WX9861,WX9859,WX9857,WX9855,WX9853,WX9851,WX9849,WX9847
	,WX9845,WX9843,WX9841,WX9839,WX9837,WX9835,WX9833,WX9831
	,WX9829,WX9827,WX9825,WX9823,WX9821,WX9819,WX9817,WX9815
	,WX9813,WX9811,WX9809,WX9807,WX9805,WX9803,WX9801,WX9799
	,WX9797,WX9795,WX9793,WX9791,WX9789,WX9787,WX9785,WX9783
	,WX9781,WX9779,WX9777,WX9775,WX9773,WX9771,WX9769,WX9767
	,WX9765,WX9763,WX9761,WX9759,WX9595,WX9593,WX9591,WX9589
	,WX9587,WX9585,WX9583,WX9581,WX9579,WX9577,WX9575,WX9573
	,WX9571,WX9569,WX9567,WX9565,WX9563,WX9561,WX9559,WX9557
	,WX9555,WX9553,WX9551,WX9549,WX9547,WX9545,WX9543,WX9541
	,WX9539,WX9537,WX9535,WX8656,WX8654,WX8652,WX8650,WX8648
	,WX8646,WX8644,WX8642,WX8640,WX8638,WX8636,WX8634,WX8632
	,WX8630,WX8628,WX8626,WX8624,WX8622,WX8620,WX8618,WX8616
	,WX8614,WX8612,WX8610,WX8608,WX8606,WX8604,WX8602,WX8600
	,WX8598,WX8596,WX8594,WX8592,WX8590,WX8588,WX8586,WX8584
	,WX8582,WX8580,WX8578,WX8576,WX8574,WX8572,WX8570,WX8568
	,WX8566,WX8564,WX8562,WX8560,WX8558,WX8556,WX8554,WX8552
	,WX8550,WX8548,WX8546,WX8544,WX8542,WX8540,WX8538,WX8536
	,WX8534,WX8532,WX8530,WX8528,WX8526,WX8524,WX8522,WX8520
	,WX8518,WX8516,WX8514,WX8512,WX8510,WX8508,WX8506,WX8504
	,WX8502,WX8500,WX8498,WX8496,WX8494,WX8492,WX8490,WX8488
	,WX8486,WX8484,WX8482,WX8480,WX8478,WX8476,WX8474,WX8472
	,WX8470,WX8468,WX8466,WX8302,WX8300,WX8298,WX8296,WX8294
	,WX8292,WX8290,WX8288,WX8286,WX8284,WX8282,WX8280,WX8278
	,WX8276,WX8274,WX8272,WX8270,WX8268,WX8266,WX8264,WX8262
	,WX8260,WX8258,WX8256,WX8254,WX8252,WX8250,WX8248,WX8246
	,WX8244,WX8242,WX7363,WX7361,WX7359,WX7357,WX7355,WX7353
	,WX7351,WX7349,WX7347,WX7345,WX7343,WX7341,WX7339,WX7337
	,WX7335,WX7333,WX7331,WX7329,WX7327,WX7325,WX7323,WX7321
	,WX7319,WX7317,WX7315,WX7313,WX7311,WX7309,WX7307,WX7305
	,WX7303,WX7301,WX7299,WX7297,WX7295,WX7293,WX7291,WX7289
	,WX7287,WX7285,WX7283,WX7281,WX7279,WX7277,WX7275,WX7273
	,WX7271,WX7269,WX7267,WX7265,WX7263,WX7261,WX7259,WX7257
	,WX7255,WX7253,WX7251,WX7249,WX7247,WX7245,WX7243,WX7241
	,WX7239,WX7237,WX7235,WX7233,WX7231,WX7229,WX7227,WX7225
	,WX7223,WX7221,WX7219,WX7217,WX7215,WX7213,WX7211,WX7209
	,WX7207,WX7205,WX7203,WX7201,WX7199,WX7197,WX7195,WX7193
	,WX7191,WX7189,WX7187,WX7185,WX7183,WX7181,WX7179,WX7177
	,WX7175,WX7173,WX7009,WX7007,WX7005,WX7003,WX7001,WX6999
	,WX6997,WX6995,WX6993,WX6991,WX6989,WX6987,WX6985,WX6983
	,WX6981,WX6979,WX6977,WX6975,WX6973,WX6971,WX6969,WX6967
	,WX6965,WX6963,WX6961,WX6959,WX6957,WX6955,WX6953,WX6951
	,WX6949,WX6070,WX6068,WX6066,WX6064,WX6062,WX6060,WX6058
	,WX6056,WX6054,WX6052,WX6050,WX6048,WX6046,WX6044,WX6042
	,WX6040,WX6038,WX6036,WX6034,WX6032,WX6030,WX6028,WX6026
	,WX6024,WX6022,WX6020,WX6018,WX6016,WX6014,WX6012,WX6010
	,WX6008,WX6006,WX6004,WX6002,WX6000,WX5998,WX5996,WX5994
	,WX5992,WX5990,WX5988,WX5986,WX5984,WX5982,WX5980,WX5978
	,WX5976,WX5974,WX5972,WX5970,WX5968,WX5966,WX5964,WX5962
	,WX5960,WX5958,WX5956,WX5954,WX5952,WX5950,WX5948,WX5946
	,WX5944,WX5942,WX5940,WX5938,WX5936,WX5934,WX5932,WX5930
	,WX5928,WX5926,WX5924,WX5922,WX5920,WX5918,WX5916,WX5914
	,WX5912,WX5910,WX5908,WX5906,WX5904,WX5902,WX5900,WX5898
	,WX5896,WX5894,WX5892,WX5890,WX5888,WX5886,WX5884,WX5882
	,WX5880,WX5716,WX5714,WX5712,WX5710,WX5708,WX5706,WX5704
	,WX5702,WX5700,WX5698,WX5696,WX5694,WX5692,WX5690,WX5688
	,WX5686,WX5684,WX5682,WX5680,WX5678,WX5676,WX5674,WX5672
	,WX5670,WX5668,WX5666,WX5664,WX5662,WX5660,WX5658,WX5656
	,WX4777,WX4775,WX4773,WX4771,WX4769,WX4767,WX4765,WX4763
	,WX4761,WX4759,WX4757,WX4755,WX4753,WX4751,WX4749,WX4747
	,WX4745,WX4743,WX4741,WX4739,WX4737,WX4735,WX4733,WX4731
	,WX4729,WX4727,WX4725,WX4723,WX4721,WX4719,WX4717,WX4715
	,WX4713,WX4711,WX4709,WX4707,WX4705,WX4703,WX4701,WX4699
	,WX4697,WX4695,WX4693,WX4691,WX4689,WX4687,WX4685,WX4683
	,WX4681,WX4679,WX4677,WX4675,WX4673,WX4671,WX4669,WX4667
	,WX4665,WX4663,WX4661,WX4659,WX4657,WX4655,WX4653,WX4651
	,WX4649,WX4647,WX4645,WX4643,WX4641,WX4639,WX4637,WX4635
	,WX4633,WX4631,WX4629,WX4627,WX4625,WX4623,WX4621,WX4619
	,WX4617,WX4615,WX4613,WX4611,WX4609,WX4607,WX4605,WX4603
	,WX4601,WX4599,WX4597,WX4595,WX4593,WX4591,WX4589,WX4587
	,WX4423,WX4421,WX4419,WX4417,WX4415,WX4413,WX4411,WX4409
	,WX4407,WX4405,WX4403,WX4401,WX4399,WX4397,WX4395,WX4393
	,WX4391,WX4389,WX4387,WX4385,WX4383,WX4381,WX4379,WX4377
	,WX4375,WX4373,WX4371,WX4369,WX4367,WX4365,WX4363,WX3484
	,WX3482,WX3480,WX3478,WX3476,WX3474,WX3472,WX3470,WX3468
	,WX3466,WX3464,WX3462,WX3460,WX3458,WX3456,WX3454,WX3452
	,WX3450,WX3448,WX3446,WX3444,WX3442,WX3440,WX3438,WX3436
	,WX3434,WX3432,WX3430,WX3428,WX3426,WX3424,WX3422,WX3420
	,WX3418,WX3416,WX3414,WX3412,WX3410,WX3408,WX3406,WX3404
	,WX3402,WX3400,WX3398,WX3396,WX3394,WX3392,WX3390,WX3388
	,WX3386,WX3384,WX3382,WX3380,WX3378,WX3376,WX3374,WX3372
	,WX3370,WX3368,WX3366,WX3364,WX3362,WX3360,WX3358,WX3356
	,WX3354,WX3352,WX3350,WX3348,WX3346,WX3344,WX3342,WX3340
	,WX3338,WX3336,WX3334,WX3332,WX3330,WX3328,WX3326,WX3324
	,WX3322,WX3320,WX3318,WX3316,WX3314,WX3312,WX3310,WX3308
	,WX3306,WX3304,WX3302,WX3300,WX3298,WX3296,WX3294,WX3130
	,WX3128,WX3126,WX3124,WX3122,WX3120,WX3118,WX3116,WX3114
	,WX3112,WX3110,WX3108,WX3106,WX3104,WX3102,WX3100,WX3098
	,WX3096,WX3094,WX3092,WX3090,WX3088,WX3086,WX3084,WX3082
	,WX3080,WX3078,WX3076,WX3074,WX3072,WX3070,WX2191,WX2189
	,WX2187,WX2185,WX2183,WX2181,WX2179,WX2177,WX2175,WX2173
	,WX2171,WX2169,WX2167,WX2165,WX2163,WX2161,WX2159,WX2157
	,WX2155,WX2153,WX2151,WX2149,WX2147,WX2145,WX2143,WX2141
	,WX2139,WX2137,WX2135,WX2133,WX2131,WX2129,WX2127,WX2125
	,WX2123,WX2121,WX2119,WX2117,WX2115,WX2113,WX2111,WX2109
	,WX2107,WX2105,WX2103,WX2101,WX2099,WX2097,WX2095,WX2093
	,WX2091,WX2089,WX2087,WX2085,WX2083,WX2081,WX2079,WX2077
	,WX2075,WX2073,WX2071,WX2069,WX2067,WX2065,WX2063,WX2061
	,WX2059,WX2057,WX2055,WX2053,WX2051,WX2049,WX2047,WX2045
	,WX2043,WX2041,WX2039,WX2037,WX2035,WX2033,WX2031,WX2029
	,WX2027,WX2025,WX2023,WX2021,WX2019,WX2017,WX2015,WX2013
	,WX2011,WX2009,WX2007,WX2005,WX2003,WX2001,WX1837,WX1835
	,WX1833,WX1831,WX1829,WX1827,WX1825,WX1823,WX1821,WX1819
	,WX1817,WX1815,WX1813,WX1811,WX1809,WX1807,WX1805,WX1803
	,WX1801,WX1799,WX1797,WX1795,WX1793,WX1791,WX1789,WX1787
	,WX1785,WX1783,WX1781,WX1779,WX1777,WX898,WX896,WX894
	,WX892,WX890,WX888,WX886,WX884,WX882,WX880,WX878
	,WX876,WX874,WX872,WX870,WX868,WX866,WX864,WX862
	,WX860,WX858,WX856,WX854,WX852,WX850,WX848,WX846
	,WX844,WX842,WX840,WX838,WX836,WX834,WX832,WX830
	,WX828,WX826,WX824,WX822,WX820,WX818,WX816,WX814
	,WX812,WX810,WX808,WX806,WX804,WX802,WX800,WX798
	,WX796,WX794,WX792,WX790,WX788,WX786,WX784,WX782
	,WX780,WX778,WX776,WX774,WX772,WX770,WX768,WX766
	,WX764,WX762,WX760,WX758,WX756,WX754,WX752,WX750
	,WX748,WX746,WX744,WX742,WX740,WX738,WX736,WX734
	,WX732,WX730,WX728,WX726,WX724,WX722,WX720,WX718
	,WX716,WX714,WX712,WX710,WX708,WX544,WX542,WX540
	,WX538,WX536,WX534,WX532,WX530,WX528,WX526,WX524
	,WX522,WX520,WX518,WX516,WX514,WX512,WX510,WX508
	,WX506,WX504,WX502,WX500,WX498,WX496,WX494,WX492
	,WX490,WX488,WX486,WX484,WX483,II2003,II2034,II2065
	,II2096,II2127,II2158,II2189,II2220,II2251,II2282,II2313
	,II2344,II2375,II2406,II2437,II2468,II2499,II2530,II2561
	,II2592,II2623,II2654,II2685,II2716,II2747,II2778,II2809
	,II2840,II2871,II2902,II2933,II2964,WX612,WX613,WX614
	,WX615,WX616,WX617,WX618,WX619,WX620,WX621,WX622
	,WX623,WX624,WX625,WX626,WX627,WX628,WX629,WX630
	,WX631,WX632,WX633,WX634,WX635,WX636,WX637,WX638
	,WX639,WX640,WX641,WX642,WX643,WX1776,II6008,II6039
	,II6070,II6101,II6132,II6163,II6194,II6225,II6256,II6287
	,II6318,II6349,II6380,II6411,II6442,II6473,II6504,II6535
	,II6566,II6597,II6628,II6659,II6690,II6721,II6752,II6783
	,II6814,II6845,II6876,II6907,II6938,II6969,WX1905,WX1906
	,WX1907,WX1908,WX1909,WX1910,WX1911,WX1912,WX1913,WX1914
	,WX1915,WX1916,WX1917,WX1918,WX1919,WX1920,WX1921,WX1922
	,WX1923,WX1924,WX1925,WX1926,WX1927,WX1928,WX1929,WX1930
	,WX1931,WX1932,WX1933,WX1934,WX1935,WX1936,WX3069,II10013
	,II10044,II10075,II10106,II10137,II10168,II10199,II10230,II10261
	,II10292,II10323,II10354,II10385,II10416,II10447,II10478,II10509
	,II10540,II10571,II10602,II10633,II10664,II10695,II10726,II10757
	,II10788,II10819,II10850,II10881,II10912,II10943,II10974,WX3198
	,WX3199,WX3200,WX3201,WX3202,WX3203,WX3204,WX3205,WX3206
	,WX3207,WX3208,WX3209,WX3210,WX3211,WX3212,WX3213,WX3214
	,WX3215,WX3216,WX3217,WX3218,WX3219,WX3220,WX3221,WX3222
	,WX3223,WX3224,WX3225,WX3226,WX3227,WX3228,WX3229,WX4362
	,II14018,II14049,II14080,II14111,II14142,II14173,II14204,II14235
	,II14266,II14297,II14328,II14359,II14390,II14421,II14452,II14483
	,II14514,II14545,II14576,II14607,II14638,II14669,II14700,II14731
	,II14762,II14793,II14824,II14855,II14886,II14917,II14948,II14979
	,WX4491,WX4492,WX4493,WX4494,WX4495,WX4496,WX4497,WX4498
	,WX4499,WX4500,WX4501,WX4502,WX4503,WX4504,WX4505,WX4506
	,WX4507,WX4508,WX4509,WX4510,WX4511,WX4512,WX4513,WX4514
	,WX4515,WX4516,WX4517,WX4518,WX4519,WX4520,WX4521,WX4522
	,WX5655,II18023,II18054,II18085,II18116,II18147,II18178,II18209
	,II18240,II18271,II18302,II18333,II18364,II18395,II18426,II18457
	,II18488,II18519,II18550,II18581,II18612,II18643,II18674,II18705
	,II18736,II18767,II18798,II18829,II18860,II18891,II18922,II18953
	,II18984,WX5784,WX5785,WX5786,WX5787,WX5788,WX5789,WX5790
	,WX5791,WX5792,WX5793,WX5794,WX5795,WX5796,WX5797,WX5798
	,WX5799,WX5800,WX5801,WX5802,WX5803,WX5804,WX5805,WX5806
	,WX5807,WX5808,WX5809,WX5810,WX5811,WX5812,WX5813,WX5814
	,WX5815,WX6948,II22028,II22059,II22090,II22121,II22152,II22183
	,II22214,II22245,II22276,II22307,II22338,II22369,II22400,II22431
	,II22462,II22493,II22524,II22555,II22586,II22617,II22648,II22679
	,II22710,II22741,II22772,II22803,II22834,II22865,II22896,II22927
	,II22958,II22989,WX7077,WX7078,WX7079,WX7080,WX7081,WX7082
	,WX7083,WX7084,WX7085,WX7086,WX7087,WX7088,WX7089,WX7090
	,WX7091,WX7092,WX7093,WX7094,WX7095,WX7096,WX7097,WX7098
	,WX7099,WX7100,WX7101,WX7102,WX7103,WX7104,WX7105,WX7106
	,WX7107,WX7108,WX8241,II26033,II26064,II26095,II26126,II26157
	,II26188,II26219,II26250,II26281,II26312,II26343,II26374,II26405
	,II26436,II26467,II26498,II26529,II26560,II26591,II26622,II26653
	,II26684,II26715,II26746,II26777,II26808,II26839,II26870,II26901
	,II26932,II26963,II26994,WX8370,WX8371,WX8372,WX8373,WX8374
	,WX8375,WX8376,WX8377,WX8378,WX8379,WX8380,WX8381,WX8382
	,WX8383,WX8384,WX8385,WX8386,WX8387,WX8388,WX8389,WX8390
	,WX8391,WX8392,WX8393,WX8394,WX8395,WX8396,WX8397,WX8398
	,WX8399,WX8400,WX8401,WX9534,II30038,II30069,II30100,II30131
	,II30162,II30193,II30224,II30255,II30286,II30317,II30348,II30379
	,II30410,II30441,II30472,II30503,II30534,II30565,II30596,II30627
	,II30658,II30689,II30720,II30751,II30782,II30813,II30844,II30875
	,II30906,II30937,II30968,II30999,WX9663,WX9664,WX9665,WX9666
	,WX9667,WX9668,WX9669,WX9670,WX9671,WX9672,WX9673,WX9674
	,WX9675,WX9676,WX9677,WX9678,WX9679,WX9680,WX9681,WX9682
	,WX9683,WX9684,WX9685,WX9686,WX9687,WX9688,WX9689,WX9690
	,WX9691,WX9692,WX9693,WX9694,WX10827,II34043,II34074,II34105
	,II34136,II34167,II34198,II34229,II34260,II34291,II34322,II34353
	,II34384,II34415,II34446,II34477,II34508,II34539,II34570,II34601
	,II34632,II34663,II34694,II34725,II34756,II34787,II34818,II34849
	,II34880,II34911,II34942,II34973,II35004,WX10956,WX10957,WX10958
	,WX10959,WX10960,WX10961,WX10962,WX10963,WX10964,WX10965,WX10966
	,WX10967,WX10968,WX10969,WX10970,WX10971,WX10972,WX10973,WX10974
	,WX10975,WX10976,WX10977,WX10978,WX10979,WX10980,WX10981,WX10982
	,WX10983,WX10984,WX10985,WX10986,WX10987,WX10815,WX10801,WX10787
	,WX10773,WX10759,WX10745,WX10731,WX10717,WX10703,WX10689,WX10675
	,WX10661,WX10647,WX10633,WX10619,WX10605,WX10591,WX10577,WX10563
	,WX10549,WX10535,WX10521,WX10507,WX10493,WX10479,WX10465,WX10451
	,WX10437,WX10423,WX10409,WX10395,WX10381,WX9522,WX9508,WX9494
	,WX9480,WX9466,WX9452,WX9438,WX9424,WX9410,WX9396,WX9382
	,WX9368,WX9354,WX9340,WX9326,WX9312,WX9298,WX9284,WX9270
	,WX9256,WX9242,WX9228,WX9214,WX9200,WX9186,WX9172,WX9158
	,WX9144,WX9130,WX9116,WX9102,WX9088,WX8229,WX8215,WX8201
	,WX8187,WX8173,WX8159,WX8145,WX8131,WX8117,WX8103,WX8089
	,WX8075,WX8061,WX8047,WX8033,WX8019,WX8005,WX7991,WX7977
	,WX7963,WX7949,WX7935,WX7921,WX7907,WX7893,WX7879,WX7865
	,WX7851,WX7837,WX7823,WX7809,WX7795,WX6936,WX6922,WX6908
	,WX6894,WX6880,WX6866,WX6852,WX6838,WX6824,WX6810,WX6796
	,WX6782,WX6768,WX6754,WX6740,WX6726,WX6712,WX6698,WX6684
	,WX6670,WX6656,WX6642,WX6628,WX6614,WX6600,WX6586,WX6572
	,WX6558,WX6544,WX6530,WX6516,WX6502,WX5643,WX5629,WX5615
	,WX5601,WX5587,WX5573,WX5559,WX5545,WX5531,WX5517,WX5503
	,WX5489,WX5475,WX5461,WX5447,WX5433,WX5419,WX5405,WX5391
	,WX5377,WX5363,WX5349,WX5335,WX5321,WX5307,WX5293,WX5279
	,WX5265,WX5251,WX5237,WX5223,WX5209,WX4350,WX4336,WX4322
	,WX4308,WX4294,WX4280,WX4266,WX4252,WX4238,WX4224,WX4210
	,WX4196,WX4182,WX4168,WX4154,WX4140,WX4126,WX4112,WX4098
	,WX4084,WX4070,WX4056,WX4042,WX4028,WX4014,WX4000,WX3986
	,WX3972,WX3958,WX3944,WX3930,WX3916,WX3057,WX3043,WX3029
	,WX3015,WX3001,WX2987,WX2973,WX2959,WX2945,WX2931,WX2917
	,WX2903,WX2889,WX2875,WX2861,WX2847,WX2833,WX2819,WX2805
	,WX2791,WX2777,WX2763,WX2749,WX2735,WX2721,WX2707,WX2693
	,WX2679,WX2665,WX2651,WX2637,WX2623,WX1764,WX1750,WX1736
	,WX1722,WX1708,WX1694,WX1680,WX1666,WX1652,WX1638,WX1624
	,WX1610,WX1596,WX1582,WX1568,WX1554,WX1540,WX1526,WX1512
	,WX1498,WX1484,WX1470,WX1456,WX1442,WX1428,WX1414,WX1400
	,WX1386,WX1372,WX1358,WX1344,WX1330,WX471,WX457,WX443
	,WX429,WX415,WX401,WX387,WX373,WX359,WX345,WX331
	,WX317,WX303,WX289,WX275,WX261,WX247,WX233,WX219
	,WX205,WX191,WX177,WX163,WX149,WX135,WX121,WX107
	,WX93,WX79,WX65,WX51,WX37,WX10823,WX10819,WX10809
	,WX10805,WX10795,WX10791,WX10781,WX10777,WX10767,WX10763,WX10753
	,WX10749,WX10739,WX10735,WX10725,WX10721,WX10711,WX10707,WX10697
	,WX10693,WX10683,WX10679,WX10669,WX10665,WX10655,WX10651,WX10641
	,WX10637,WX10627,WX10623,WX10613,WX10609,WX10599,WX10595,WX10585
	,WX10581,WX10571,WX10567,WX10557,WX10553,WX10543,WX10539,WX10529
	,WX10525,WX10515,WX10511,WX10501,WX10497,WX10487,WX10483,WX10473
	,WX10469,WX10459,WX10455,WX10445,WX10441,WX10431,WX10427,WX10417
	,WX10413,WX10403,WX10399,WX10389,WX10385,WX11570,WX11563,WX11556
	,WX11549,WX11542,WX11535,WX11528,WX11521,WX11514,WX11507,WX11500
	,WX11493,WX11486,WX11479,WX11472,WX11465,WX11458,WX11451,WX11444
	,WX11437,WX11430,WX11423,WX11416,WX11409,WX11402,WX11395,WX11388
	,WX11381,WX11374,WX11367,WX11360,WX11353,WX9530,WX9526,WX9516
	,WX9512,WX9502,WX9498,WX9488,WX9484,WX9474,WX9470,WX9460
	,WX9456,WX9446,WX9442,WX9432,WX9428,WX9418,WX9414,WX9404
	,WX9400,WX9390,WX9386,WX9376,WX9372,WX9362,WX9358,WX9348
	,WX9344,WX9334,WX9330,WX9320,WX9316,WX9306,WX9302,WX9292
	,WX9288,WX9278,WX9274,WX9264,WX9260,WX9250,WX9246,WX9236
	,WX9232,WX9222,WX9218,WX9208,WX9204,WX9194,WX9190,WX9180
	,WX9176,WX9166,WX9162,WX9152,WX9148,WX9138,WX9134,WX9124
	,WX9120,WX9110,WX9106,WX9096,WX9092,WX10277,WX10270,WX10263
	,WX10256,WX10249,WX10242,WX10235,WX10228,WX10221,WX10214,WX10207
	,WX10200,WX10193,WX10186,WX10179,WX10172,WX10165,WX10158,WX10151
	,WX10144,WX10137,WX10130,WX10123,WX10116,WX10109,WX10102,WX10095
	,WX10088,WX10081,WX10074,WX10067,WX10060,WX8237,WX8233,WX8223
	,WX8219,WX8209,WX8205,WX8195,WX8191,WX8181,WX8177,WX8167
	,WX8163,WX8153,WX8149,WX8139,WX8135,WX8125,WX8121,WX8111
	,WX8107,WX8097,WX8093,WX8083,WX8079,WX8069,WX8065,WX8055
	,WX8051,WX8041,WX8037,WX8027,WX8023,WX8013,WX8009,WX7999
	,WX7995,WX7985,WX7981,WX7971,WX7967,WX7957,WX7953,WX7943
	,WX7939,WX7929,WX7925,WX7915,WX7911,WX7901,WX7897,WX7887
	,WX7883,WX7873,WX7869,WX7859,WX7855,WX7845,WX7841,WX7831
	,WX7827,WX7817,WX7813,WX7803,WX7799,WX8984,WX8977,WX8970
	,WX8963,WX8956,WX8949,WX8942,WX8935,WX8928,WX8921,WX8914
	,WX8907,WX8900,WX8893,WX8886,WX8879,WX8872,WX8865,WX8858
	,WX8851,WX8844,WX8837,WX8830,WX8823,WX8816,WX8809,WX8802
	,WX8795,WX8788,WX8781,WX8774,WX8767,WX6944,WX6940,WX6930
	,WX6926,WX6916,WX6912,WX6902,WX6898,WX6888,WX6884,WX6874
	,WX6870,WX6860,WX6856,WX6846,WX6842,WX6832,WX6828,WX6818
	,WX6814,WX6804,WX6800,WX6790,WX6786,WX6776,WX6772,WX6762
	,WX6758,WX6748,WX6744,WX6734,WX6730,WX6720,WX6716,WX6706
	,WX6702,WX6692,WX6688,WX6678,WX6674,WX6664,WX6660,WX6650
	,WX6646,WX6636,WX6632,WX6622,WX6618,WX6608,WX6604,WX6594
	,WX6590,WX6580,WX6576,WX6566,WX6562,WX6552,WX6548,WX6538
	,WX6534,WX6524,WX6520,WX6510,WX6506,WX7691,WX7684,WX7677
	,WX7670,WX7663,WX7656,WX7649,WX7642,WX7635,WX7628,WX7621
	,WX7614,WX7607,WX7600,WX7593,WX7586,WX7579,WX7572,WX7565
	,WX7558,WX7551,WX7544,WX7537,WX7530,WX7523,WX7516,WX7509
	,WX7502,WX7495,WX7488,WX7481,WX7474,WX5651,WX5647,WX5637
	,WX5633,WX5623,WX5619,WX5609,WX5605,WX5595,WX5591,WX5581
	,WX5577,WX5567,WX5563,WX5553,WX5549,WX5539,WX5535,WX5525
	,WX5521,WX5511,WX5507,WX5497,WX5493,WX5483,WX5479,WX5469
	,WX5465,WX5455,WX5451,WX5441,WX5437,WX5427,WX5423,WX5413
	,WX5409,WX5399,WX5395,WX5385,WX5381,WX5371,WX5367,WX5357
	,WX5353,WX5343,WX5339,WX5329,WX5325,WX5315,WX5311,WX5301
	,WX5297,WX5287,WX5283,WX5273,WX5269,WX5259,WX5255,WX5245
	,WX5241,WX5231,WX5227,WX5217,WX5213,WX6398,WX6391,WX6384
	,WX6377,WX6370,WX6363,WX6356,WX6349,WX6342,WX6335,WX6328
	,WX6321,WX6314,WX6307,WX6300,WX6293,WX6286,WX6279,WX6272
	,WX6265,WX6258,WX6251,WX6244,WX6237,WX6230,WX6223,WX6216
	,WX6209,WX6202,WX6195,WX6188,WX6181,WX4358,WX4354,WX4344
	,WX4340,WX4330,WX4326,WX4316,WX4312,WX4302,WX4298,WX4288
	,WX4284,WX4274,WX4270,WX4260,WX4256,WX4246,WX4242,WX4232
	,WX4228,WX4218,WX4214,WX4204,WX4200,WX4190,WX4186,WX4176
	,WX4172,WX4162,WX4158,WX4148,WX4144,WX4134,WX4130,WX4120
	,WX4116,WX4106,WX4102,WX4092,WX4088,WX4078,WX4074,WX4064
	,WX4060,WX4050,WX4046,WX4036,WX4032,WX4022,WX4018,WX4008
	,WX4004,WX3994,WX3990,WX3980,WX3976,WX3966,WX3962,WX3952
	,WX3948,WX3938,WX3934,WX3924,WX3920,WX5105,WX5098,WX5091
	,WX5084,WX5077,WX5070,WX5063,WX5056,WX5049,WX5042,WX5035
	,WX5028,WX5021,WX5014,WX5007,WX5000,WX4993,WX4986,WX4979
	,WX4972,WX4965,WX4958,WX4951,WX4944,WX4937,WX4930,WX4923
	,WX4916,WX4909,WX4902,WX4895,WX4888,WX3065,WX3061,WX3051
	,WX3047,WX3037,WX3033,WX3023,WX3019,WX3009,WX3005,WX2995
	,WX2991,WX2981,WX2977,WX2967,WX2963,WX2953,WX2949,WX2939
	,WX2935,WX2925,WX2921,WX2911,WX2907,WX2897,WX2893,WX2883
	,WX2879,WX2869,WX2865,WX2855,WX2851,WX2841,WX2837,WX2827
	,WX2823,WX2813,WX2809,WX2799,WX2795,WX2785,WX2781,WX2771
	,WX2767,WX2757,WX2753,WX2743,WX2739,WX2729,WX2725,WX2715
	,WX2711,WX2701,WX2697,WX2687,WX2683,WX2673,WX2669,WX2659
	,WX2655,WX2645,WX2641,WX2631,WX2627,WX3812,WX3805,WX3798
	,WX3791,WX3784,WX3777,WX3770,WX3763,WX3756,WX3749,WX3742
	,WX3735,WX3728,WX3721,WX3714,WX3707,WX3700,WX3693,WX3686
	,WX3679,WX3672,WX3665,WX3658,WX3651,WX3644,WX3637,WX3630
	,WX3623,WX3616,WX3609,WX3602,WX3595,WX1772,WX1768,WX1758
	,WX1754,WX1744,WX1740,WX1730,WX1726,WX1716,WX1712,WX1702
	,WX1698,WX1688,WX1684,WX1674,WX1670,WX1660,WX1656,WX1646
	,WX1642,WX1632,WX1628,WX1618,WX1614,WX1604,WX1600,WX1590
	,WX1586,WX1576,WX1572,WX1562,WX1558,WX1548,WX1544,WX1534
	,WX1530,WX1520,WX1516,WX1506,WX1502,WX1492,WX1488,WX1478
	,WX1474,WX1464,WX1460,WX1450,WX1446,WX1436,WX1432,WX1422
	,WX1418,WX1408,WX1404,WX1394,WX1390,WX1380,WX1376,WX1366
	,WX1362,WX1352,WX1348,WX1338,WX1334,WX2519,WX2512,WX2505
	,WX2498,WX2491,WX2484,WX2477,WX2470,WX2463,WX2456,WX2449
	,WX2442,WX2435,WX2428,WX2421,WX2414,WX2407,WX2400,WX2393
	,WX2386,WX2379,WX2372,WX2365,WX2358,WX2351,WX2344,WX2337
	,WX2330,WX2323,WX2316,WX2309,WX2302,WX479,WX475,WX465
	,WX461,WX451,WX447,WX437,WX433,WX423,WX419,WX409
	,WX405,WX395,WX391,WX381,WX377,WX367,WX363,WX353
	,WX349,WX339,WX335,WX325,WX321,WX311,WX307,WX297
	,WX293,WX283,WX279,WX269,WX265,WX255,WX251,WX241
	,WX237,WX227,WX223,WX213,WX209,WX199,WX195,WX185
	,WX181,WX171,WX167,WX157,WX153,WX143,WX139,WX129
	,WX125,WX115,WX111,WX101,WX97,WX87,WX83,WX73
	,WX69,WX59,WX55,WX45,WX41,WX1226,WX1219,WX1212
	,WX1205,WX1198,WX1191,WX1184,WX1177,WX1170,WX1163,WX1156
	,WX1149,WX1142,WX1135,WX1128,WX1121,WX1114,WX1107,WX1100
	,WX1093,WX1086,WX1079,WX1072,WX1065,WX1058,WX1051,WX1044
	,WX1037,WX1030,WX1023,WX1016,WX1009,II35006,II34975,II34944
	,II34913,II34882,II34851,II34820,II34789,II34758,II34727,II34696
	,II34665,II34634,II34603,II34572,II34541,II34510,II34479,II34448
	,II34417,II34386,II34355,II34324,II34293,II34262,II34231,II34200
	,II34169,II34138,II34107,II34076,II34045,II34989,II34958,II34927
	,II34896,II34865,II34834,II34803,II34772,II34741,II34710,II34679
	,II34648,II34617,II34586,II34555,II34524,II34493,II34462,II34431
	,II34400,II34369,II34338,II34307,II34276,II34245,II34214,II34183
	,II34152,II34121,II34090,II34059,II34028,WX10821,WX10807,WX10793
	,WX10779,WX10765,WX10751,WX10737,WX10723,WX10709,WX10695,WX10681
	,WX10667,WX10653,WX10639,WX10625,WX10611,WX10597,WX10583,WX10569
	,WX10555,WX10541,WX10527,WX10513,WX10499,WX10485,WX10471,WX10457
	,WX10443,WX10429,WX10415,WX10401,WX10387,II31001,II30970,II30939
	,II30908,II30877,II30846,II30815,II30784,II30753,II30722,II30691
	,II30660,II30629,II30598,II30567,II30536,II30505,II30474,II30443
	,II30412,II30381,II30350,II30319,II30288,II30257,II30226,II30195
	,II30164,II30133,II30102,II30071,II30040,II30984,II30953,II30922
	,II30891,II30860,II30829,II30798,II30767,II30736,II30705,II30674
	,II30643,II30612,II30581,II30550,II30519,II30488,II30457,II30426
	,II30395,II30364,II30333,II30302,II30271,II30240,II30209,II30178
	,II30147,II30116,II30085,II30054,II30023,WX9528,WX9514,WX9500
	,WX9486,WX9472,WX9458,WX9444,WX9430,WX9416,WX9402,WX9388
	,WX9374,WX9360,WX9346,WX9332,WX9318,WX9304,WX9290,WX9276
	,WX9262,WX9248,WX9234,WX9220,WX9206,WX9192,WX9178,WX9164
	,WX9150,WX9136,WX9122,WX9108,WX9094,II26996,II26965,II26934
	,II26903,II26872,II26841,II26810,II26779,II26748,II26717,II26686
	,II26655,II26624,II26593,II26562,II26531,II26500,II26469,II26438
	,II26407,II26376,II26345,II26314,II26283,II26252,II26221,II26190
	,II26159,II26128,II26097,II26066,II26035,II26979,II26948,II26917
	,II26886,II26855,II26824,II26793,II26762,II26731,II26700,II26669
	,II26638,II26607,II26576,II26545,II26514,II26483,II26452,II26421
	,II26390,II26359,II26328,II26297,II26266,II26235,II26204,II26173
	,II26142,II26111,II26080,II26049,II26018,WX8235,WX8221,WX8207
	,WX8193,WX8179,WX8165,WX8151,WX8137,WX8123,WX8109,WX8095
	,WX8081,WX8067,WX8053,WX8039,WX8025,WX8011,WX7997,WX7983
	,WX7969,WX7955,WX7941,WX7927,WX7913,WX7899,WX7885,WX7871
	,WX7857,WX7843,WX7829,WX7815,WX7801,II22991,II22960,II22929
	,II22898,II22867,II22836,II22805,II22774,II22743,II22712,II22681
	,II22650,II22619,II22588,II22557,II22526,II22495,II22464,II22433
	,II22402,II22371,II22340,II22309,II22278,II22247,II22216,II22185
	,II22154,II22123,II22092,II22061,II22030,II22974,II22943,II22912
	,II22881,II22850,II22819,II22788,II22757,II22726,II22695,II22664
	,II22633,II22602,II22571,II22540,II22509,II22478,II22447,II22416
	,II22385,II22354,II22323,II22292,II22261,II22230,II22199,II22168
	,II22137,II22106,II22075,II22044,II22013,WX6942,WX6928,WX6914
	,WX6900,WX6886,WX6872,WX6858,WX6844,WX6830,WX6816,WX6802
	,WX6788,WX6774,WX6760,WX6746,WX6732,WX6718,WX6704,WX6690
	,WX6676,WX6662,WX6648,WX6634,WX6620,WX6606,WX6592,WX6578
	,WX6564,WX6550,WX6536,WX6522,WX6508,II18986,II18955,II18924
	,II18893,II18862,II18831,II18800,II18769,II18738,II18707,II18676
	,II18645,II18614,II18583,II18552,II18521,II18490,II18459,II18428
	,II18397,II18366,II18335,II18304,II18273,II18242,II18211,II18180
	,II18149,II18118,II18087,II18056,II18025,II18969,II18938,II18907
	,II18876,II18845,II18814,II18783,II18752,II18721,II18690,II18659
	,II18628,II18597,II18566,II18535,II18504,II18473,II18442,II18411
	,II18380,II18349,II18318,II18287,II18256,II18225,II18194,II18163
	,II18132,II18101,II18070,II18039,II18008,WX5649,WX5635,WX5621
	,WX5607,WX5593,WX5579,WX5565,WX5551,WX5537,WX5523,WX5509
	,WX5495,WX5481,WX5467,WX5453,WX5439,WX5425,WX5411,WX5397
	,WX5383,WX5369,WX5355,WX5341,WX5327,WX5313,WX5299,WX5285
	,WX5271,WX5257,WX5243,WX5229,WX5215,II14981,II14950,II14919
	,II14888,II14857,II14826,II14795,II14764,II14733,II14702,II14671
	,II14640,II14609,II14578,II14547,II14516,II14485,II14454,II14423
	,II14392,II14361,II14330,II14299,II14268,II14237,II14206,II14175
	,II14144,II14113,II14082,II14051,II14020,II14964,II14933,II14902
	,II14871,II14840,II14809,II14778,II14747,II14716,II14685,II14654
	,II14623,II14592,II14561,II14530,II14499,II14468,II14437,II14406
	,II14375,II14344,II14313,II14282,II14251,II14220,II14189,II14158
	,II14127,II14096,II14065,II14034,II14003,WX4356,WX4342,WX4328
	,WX4314,WX4300,WX4286,WX4272,WX4258,WX4244,WX4230,WX4216
	,WX4202,WX4188,WX4174,WX4160,WX4146,WX4132,WX4118,WX4104
	,WX4090,WX4076,WX4062,WX4048,WX4034,WX4020,WX4006,WX3992
	,WX3978,WX3964,WX3950,WX3936,WX3922,II10976,II10945,II10914
	,II10883,II10852,II10821,II10790,II10759,II10728,II10697,II10666
	,II10635,II10604,II10573,II10542,II10511,II10480,II10449,II10418
	,II10387,II10356,II10325,II10294,II10263,II10232,II10201,II10170
	,II10139,II10108,II10077,II10046,II10015,II10959,II10928,II10897
	,II10866,II10835,II10804,II10773,II10742,II10711,II10680,II10649
	,II10618,II10587,II10556,II10525,II10494,II10463,II10432,II10401
	,II10370,II10339,II10308,II10277,II10246,II10215,II10184,II10153
	,II10122,II10091,II10060,II10029,II9998,WX3063,WX3049,WX3035
	,WX3021,WX3007,WX2993,WX2979,WX2965,WX2951,WX2937,WX2923
	,WX2909,WX2895,WX2881,WX2867,WX2853,WX2839,WX2825,WX2811
	,WX2797,WX2783,WX2769,WX2755,WX2741,WX2727,WX2713,WX2699
	,WX2685,WX2671,WX2657,WX2643,WX2629,II6971,II6940,II6909
	,II6878,II6847,II6816,II6785,II6754,II6723,II6692,II6661
	,II6630,II6599,II6568,II6537,II6506,II6475,II6444,II6413
	,II6382,II6351,II6320,II6289,II6258,II6227,II6196,II6165
	,II6134,II6103,II6072,II6041,II6010,II6954,II6923,II6892
	,II6861,II6830,II6799,II6768,II6737,II6706,II6675,II6644
	,II6613,II6582,II6551,II6520,II6489,II6458,II6427,II6396
	,II6365,II6334,II6303,II6272,II6241,II6210,II6179,II6148
	,II6117,II6086,II6055,II6024,II5993,WX1770,WX1756,WX1742
	,WX1728,WX1714,WX1700,WX1686,WX1672,WX1658,WX1644,WX1630
	,WX1616,WX1602,WX1588,WX1574,WX1560,WX1546,WX1532,WX1518
	,WX1504,WX1490,WX1476,WX1462,WX1448,WX1434,WX1420,WX1406
	,WX1392,WX1378,WX1364,WX1350,WX1336,II2966,II2935,II2904
	,II2873,II2842,II2811,II2780,II2749,II2718,II2687,II2656
	,II2625,II2594,II2563,II2532,II2501,II2470,II2439,II2408
	,II2377,II2346,II2315,II2284,II2253,II2222,II2191,II2160
	,II2129,II2098,II2067,II2036,II2005,II2949,II2918,II2887
	,II2856,II2825,II2794,II2763,II2732,II2701,II2670,II2639
	,II2608,II2577,II2546,II2515,II2484,II2453,II2422,II2391
	,II2360,II2329,II2298,II2267,II2236,II2205,II2174,II2143
	,II2112,II2081,II2050,II2019,II1988,WX477,WX463,WX449
	,WX435,WX421,WX407,WX393,WX379,WX365,WX351,WX337
	,WX323,WX309,WX295,WX281,WX267,WX253,WX239,WX225
	,WX211,WX197,WX183,WX169,WX155,WX141,WX127,WX113
	,WX99,WX85,WX71,WX57,WX43,WX10383,WX10397,WX10411
	,WX10425,WX10439,WX10453,WX10467,WX10481,WX10495,WX10509,WX10523
	,WX10537,WX10551,WX10565,WX10579,WX10593,WX10607,WX10621,WX10635
	,WX10649,WX10663,WX10677,WX10691,WX10705,WX10719,WX10733,WX10747
	,WX10761,WX10775,WX10789,WX10803,WX10817,WX9090,WX9104,WX9118
	,WX9132,WX9146,WX9160,WX9174,WX9188,WX9202,WX9216,WX9230
	,WX9244,WX9258,WX9272,WX9286,WX9300,WX9314,WX9328,WX9342
	,WX9356,WX9370,WX9384,WX9398,WX9412,WX9426,WX9440,WX9454
	,WX9468,WX9482,WX9496,WX9510,WX9524,WX7797,WX7811,WX7825
	,WX7839,WX7853,WX7867,WX7881,WX7895,WX7909,WX7923,WX7937
	,WX7951,WX7965,WX7979,WX7993,WX8007,WX8021,WX8035,WX8049
	,WX8063,WX8077,WX8091,WX8105,WX8119,WX8133,WX8147,WX8161
	,WX8175,WX8189,WX8203,WX8217,WX8231,WX6504,WX6518,WX6532
	,WX6546,WX6560,WX6574,WX6588,WX6602,WX6616,WX6630,WX6644
	,WX6658,WX6672,WX6686,WX6700,WX6714,WX6728,WX6742,WX6756
	,WX6770,WX6784,WX6798,WX6812,WX6826,WX6840,WX6854,WX6868
	,WX6882,WX6896,WX6910,WX6924,WX6938,WX5211,WX5225,WX5239
	,WX5253,WX5267,WX5281,WX5295,WX5309,WX5323,WX5337,WX5351
	,WX5365,WX5379,WX5393,WX5407,WX5421,WX5435,WX5449,WX5463
	,WX5477,WX5491,WX5505,WX5519,WX5533,WX5547,WX5561,WX5575
	,WX5589,WX5603,WX5617,WX5631,WX5645,WX3918,WX3932,WX3946
	,WX3960,WX3974,WX3988,WX4002,WX4016,WX4030,WX4044,WX4058
	,WX4072,WX4086,WX4100,WX4114,WX4128,WX4142,WX4156,WX4170
	,WX4184,WX4198,WX4212,WX4226,WX4240,WX4254,WX4268,WX4282
	,WX4296,WX4310,WX4324,WX4338,WX4352,WX2625,WX2639,WX2653
	,WX2667,WX2681,WX2695,WX2709,WX2723,WX2737,WX2751,WX2765
	,WX2779,WX2793,WX2807,WX2821,WX2835,WX2849,WX2863,WX2877
	,WX2891,WX2905,WX2919,WX2933,WX2947,WX2961,WX2975,WX2989
	,WX3003,WX3017,WX3031,WX3045,WX3059,WX1332,WX1346,WX1360
	,WX1374,WX1388,WX1402,WX1416,WX1430,WX1444,WX1458,WX1472
	,WX1486,WX1500,WX1514,WX1528,WX1542,WX1556,WX1570,WX1584
	,WX1598,WX1612,WX1626,WX1640,WX1654,WX1668,WX1682,WX1696
	,WX1710,WX1724,WX1738,WX1752,WX1766,WX39,WX53,WX67
	,WX81,WX95,WX109,WX123,WX137,WX151,WX165,WX179
	,WX193,WX207,WX221,WX235,WX249,WX263,WX277,WX291
	,WX305,WX319,WX333,WX347,WX361,WX375,WX389,WX403
	,WX417,WX431,WX445,WX459,WX473,WX10890,WX9597,WX8304
	,WX7011,WX5718,WX4425,WX3132,WX1839,WX546,II3710,II3703
	,II3696,II3689,II3682,II3675,II3668,II3661,II3654,II3647
	,II3640,II3633,II3626,II3619,II3612,II3605,II3598,II3591
	,II3584,II3577,II3570,II3563,II3556,II3549,II3542,II3535
	,II3528,II3521,II3514,II3500,II3485,II3470,II7715,II7708
	,II7701,II7694,II7687,II7680,II7673,II7666,II7659,II7652
	,II7645,II7638,II7631,II7624,II7617,II7610,II7603,II7596
	,II7589,II7582,II7575,II7568,II7561,II7554,II7547,II7540
	,II7533,II7526,II7519,II7505,II7490,II7475,II11720,II11713
	,II11706,II11699,II11692,II11685,II11678,II11671,II11664,II11657
	,II11650,II11643,II11636,II11629,II11622,II11615,II11608,II11601
	,II11594,II11587,II11580,II11573,II11566,II11559,II11552,II11545
	,II11538,II11531,II11524,II11510,II11495,II11480,II15725,II15718
	,II15711,II15704,II15697,II15690,II15683,II15676,II15669,II15662
	,II15655,II15648,II15641,II15634,II15627,II15620,II15613,II15606
	,II15599,II15592,II15585,II15578,II15571,II15564,II15557,II15550
	,II15543,II15536,II15529,II15515,II15500,II15485,II19730,II19723
	,II19716,II19709,II19702,II19695,II19688,II19681,II19674,II19667
	,II19660,II19653,II19646,II19639,II19632,II19625,II19618,II19611
	,II19604,II19597,II19590,II19583,II19576,II19569,II19562,II19555
	,II19548,II19541,II19534,II19520,II19505,II19490,II23735,II23728
	,II23721,II23714,II23707,II23700,II23693,II23686,II23679,II23672
	,II23665,II23658,II23651,II23644,II23637,II23630,II23623,II23616
	,II23609,II23602,II23595,II23588,II23581,II23574,II23567,II23560
	,II23553,II23546,II23539,II23525,II23510,II23495,II27740,II27733
	,II27726,II27719,II27712,II27705,II27698,II27691,II27684,II27677
	,II27670,II27663,II27656,II27649,II27642,II27635,II27628,II27621
	,II27614,II27607,II27600,II27593,II27586,II27579,II27572,II27565
	,II27558,II27551,II27544,II27530,II27515,II27500,II31745,II31738
	,II31731,II31724,II31717,II31710,II31703,II31696,II31689,II31682
	,II31675,II31668,II31661,II31654,II31647,II31640,II31633,II31626
	,II31619,II31612,II31605,II31598,II31591,II31584,II31577,II31570
	,II31563,II31556,II31549,II31535,II31520,II31505,II35750,II35743
	,II35736,II35729,II35722,II35715,II35708,II35701,II35694,II35687
	,II35680,II35673,II35666,II35659,II35652,II35645,II35638,II35631
	,II35624,II35617,II35610,II35603,II35596,II35589,II35582,II35575
	,II35568,II35561,II35554,II35540,II35525,II35510,II2004,II2035
	,II2066,II2097,II2128,II2159,II2190,II2221,II2252,II2283
	,II2314,II2345,II2376,II2407,II2438,II2469,II2500,II2531
	,II2562,II2593,II2624,II2655,II2686,II2717,II2748,II2779
	,II2810,II2841,II2872,II2903,II2934,II2965,II6009,II6040
	,II6071,II6102,II6133,II6164,II6195,II6226,II6257,II6288
	,II6319,II6350,II6381,II6412,II6443,II6474,II6505,II6536
	,II6567,II6598,II6629,II6660,II6691,II6722,II6753,II6784
	,II6815,II6846,II6877,II6908,II6939,II6970,II10014,II10045
	,II10076,II10107,II10138,II10169,II10200,II10231,II10262,II10293
	,II10324,II10355,II10386,II10417,II10448,II10479,II10510,II10541
	,II10572,II10603,II10634,II10665,II10696,II10727,II10758,II10789
	,II10820,II10851,II10882,II10913,II10944,II10975,II14019,II14050
	,II14081,II14112,II14143,II14174,II14205,II14236,II14267,II14298
	,II14329,II14360,II14391,II14422,II14453,II14484,II14515,II14546
	,II14577,II14608,II14639,II14670,II14701,II14732,II14763,II14794
	,II14825,II14856,II14887,II14918,II14949,II14980,II18024,II18055
	,II18086,II18117,II18148,II18179,II18210,II18241,II18272,II18303
	,II18334,II18365,II18396,II18427,II18458,II18489,II18520,II18551
	,II18582,II18613,II18644,II18675,II18706,II18737,II18768,II18799
	,II18830,II18861,II18892,II18923,II18954,II18985,II22029,II22060
	,II22091,II22122,II22153,II22184,II22215,II22246,II22277,II22308
	,II22339,II22370,II22401,II22432,II22463,II22494,II22525,II22556
	,II22587,II22618,II22649,II22680,II22711,II22742,II22773,II22804
	,II22835,II22866,II22897,II22928,II22959,II22990,II26034,II26065
	,II26096,II26127,II26158,II26189,II26220,II26251,II26282,II26313
	,II26344,II26375,II26406,II26437,II26468,II26499,II26530,II26561
	,II26592,II26623,II26654,II26685,II26716,II26747,II26778,II26809
	,II26840,II26871,II26902,II26933,II26964,II26995,II30039,II30070
	,II30101,II30132,II30163,II30194,II30225,II30256,II30287,II30318
	,II30349,II30380,II30411,II30442,II30473,II30504,II30535,II30566
	,II30597,II30628,II30659,II30690,II30721,II30752,II30783,II30814
	,II30845,II30876,II30907,II30938,II30969,II31000,II34044,II34075
	,II34106,II34137,II34168,II34199,II34230,II34261,II34292,II34323
	,II34354,II34385,II34416,II34447,II34478,II34509,II34540,II34571
	,II34602,II34633,II34664,II34695,II34726,II34757,II34788,II34819
	,II34850,II34881,II34912,II34943,II34974,II35005,WX10384,WX10398
	,WX10412,WX10426,WX10440,WX10454,WX10468,WX10482,WX10496,WX10510
	,WX10524,WX10538,WX10552,WX10566,WX10580,WX10594,WX10608,WX10622
	,WX10636,WX10650,WX10664,WX10678,WX10692,WX10706,WX10720,WX10734
	,WX10748,WX10762,WX10776,WX10790,WX10804,WX10818,II34494,II34463
	,II34432,II34401,II34370,II34339,II34308,II34277,II34246,II34215
	,II34184,II34153,II34122,II34091,II34060,II34029,II30489,II30458
	,II30427,II30396,II30365,II30334,II30303,II30272,II30241,II30210
	,II30179,II30148,II30117,II30086,II30055,II30024,II26484,II26453
	,II26422,II26391,II26360,II26329,II26298,II26267,II26236,II26205
	,II26174,II26143,II26112,II26081,II26050,II26019,II22479,II22448
	,II22417,II22386,II22355,II22324,II22293,II22262,II22231,II22200
	,II22169,II22138,II22107,II22076,II22045,II22014,II18474,II18443
	,II18412,II18381,II18350,II18319,II18288,II18257,II18226,II18195
	,II18164,II18133,II18102,II18071,II18040,II18009,II14469,II14438
	,II14407,II14376,II14345,II14314,II14283,II14252,II14221,II14190
	,II14159,II14128,II14097,II14066,II14035,II14004,II10464,II10433
	,II10402,II10371,II10340,II10309,II10278,II10247,II10216,II10185
	,II10154,II10123,II10092,II10061,II10030,II9999,II6459,II6428
	,II6397,II6366,II6335,II6304,II6273,II6242,II6211,II6180
	,II6149,II6118,II6087,II6056,II6025,II5994,II2454,II2423
	,II2392,II2361,II2330,II2299,II2268,II2237,II2206,II2175
	,II2144,II2113,II2082,II2051,II2020,II1989,II34990,II34959
	,II34928,II34897,II34866,II34835,II34804,II34773,II34742,II34711
	,II34680,II34649,II34618,II34587,II34556,II34525,II30985,II30954
	,II30923,II30892,II30861,II30830,II30799,II30768,II30737,II30706
	,II30675,II30644,II30613,II30582,II30551,II30520,II26980,II26949
	,II26918,II26887,II26856,II26825,II26794,II26763,II26732,II26701
	,II26670,II26639,II26608,II26577,II26546,II26515,II22975,II22944
	,II22913,II22882,II22851,II22820,II22789,II22758,II22727,II22696
	,II22665,II22634,II22603,II22572,II22541,II22510,II18970,II18939
	,II18908,II18877,II18846,II18815,II18784,II18753,II18722,II18691
	,II18660,II18629,II18598,II18567,II18536,II18505,II14965,II14934
	,II14903,II14872,II14841,II14810,II14779,II14748,II14717,II14686
	,II14655,II14624,II14593,II14562,II14531,II14500,II10960,II10929
	,II10898,II10867,II10836,II10805,II10774,II10743,II10712,II10681
	,II10650,II10619,II10588,II10557,II10526,II10495,II6955,II6924
	,II6893,II6862,II6831,II6800,II6769,II6738,II6707,II6676
	,II6645,II6614,II6583,II6552,II6521,II6490,II2950,II2919
	,II2888,II2857,II2826,II2795,II2764,II2733,II2702,II2671
	,II2640,II2609,II2578,II2547,II2516,II2485,II1990,II2021
	,II2052,II2083,II2114,II2145,II2176,II2207,II2238,II2269
	,II2300,II2331,II2362,II2393,II2424,II2455,II2486,II2517
	,II2548,II2579,II2610,II2641,II2672,II2703,II2734,II2765
	,II2796,II2827,II2858,II2889,II2920,II2951,II2002,II2033
	,II2064,II2095,II2126,II2157,II2188,II2219,II2250,II2281
	,II2312,II2343,II2374,II2405,II2436,II2467,II2498,II2529
	,II2560,II2591,II2622,II2653,II2684,II2715,II2746,II2777
	,II2808,II2839,II2870,II2901,II2932,II2963,II5995,II6026
	,II6057,II6088,II6119,II6150,II6181,II6212,II6243,II6274
	,II6305,II6336,II6367,II6398,II6429,II6460,II6491,II6522
	,II6553,II6584,II6615,II6646,II6677,II6708,II6739,II6770
	,II6801,II6832,II6863,II6894,II6925,II6956,II6007,II6038
	,II6069,II6100,II6131,II6162,II6193,II6224,II6255,II6286
	,II6317,II6348,II6379,II6410,II6441,II6472,II6503,II6534
	,II6565,II6596,II6627,II6658,II6689,II6720,II6751,II6782
	,II6813,II6844,II6875,II6906,II6937,II6968,II10000,II10031
	,II10062,II10093,II10124,II10155,II10186,II10217,II10248,II10279
	,II10310,II10341,II10372,II10403,II10434,II10465,II10496,II10527
	,II10558,II10589,II10620,II10651,II10682,II10713,II10744,II10775
	,II10806,II10837,II10868,II10899,II10930,II10961,II10012,II10043
	,II10074,II10105,II10136,II10167,II10198,II10229,II10260,II10291
	,II10322,II10353,II10384,II10415,II10446,II10477,II10508,II10539
	,II10570,II10601,II10632,II10663,II10694,II10725,II10756,II10787
	,II10818,II10849,II10880,II10911,II10942,II10973,II14005,II14036
	,II14067,II14098,II14129,II14160,II14191,II14222,II14253,II14284
	,II14315,II14346,II14377,II14408,II14439,II14470,II14501,II14532
	,II14563,II14594,II14625,II14656,II14687,II14718,II14749,II14780
	,II14811,II14842,II14873,II14904,II14935,II14966,II14017,II14048
	,II14079,II14110,II14141,II14172,II14203,II14234,II14265,II14296
	,II14327,II14358,II14389,II14420,II14451,II14482,II14513,II14544
	,II14575,II14606,II14637,II14668,II14699,II14730,II14761,II14792
	,II14823,II14854,II14885,II14916,II14947,II14978,II18010,II18041
	,II18072,II18103,II18134,II18165,II18196,II18227,II18258,II18289
	,II18320,II18351,II18382,II18413,II18444,II18475,II18506,II18537
	,II18568,II18599,II18630,II18661,II18692,II18723,II18754,II18785
	,II18816,II18847,II18878,II18909,II18940,II18971,II18022,II18053
	,II18084,II18115,II18146,II18177,II18208,II18239,II18270,II18301
	,II18332,II18363,II18394,II18425,II18456,II18487,II18518,II18549
	,II18580,II18611,II18642,II18673,II18704,II18735,II18766,II18797
	,II18828,II18859,II18890,II18921,II18952,II18983,II22015,II22046
	,II22077,II22108,II22139,II22170,II22201,II22232,II22263,II22294
	,II22325,II22356,II22387,II22418,II22449,II22480,II22511,II22542
	,II22573,II22604,II22635,II22666,II22697,II22728,II22759,II22790
	,II22821,II22852,II22883,II22914,II22945,II22976,II22027,II22058
	,II22089,II22120,II22151,II22182,II22213,II22244,II22275,II22306
	,II22337,II22368,II22399,II22430,II22461,II22492,II22523,II22554
	,II22585,II22616,II22647,II22678,II22709,II22740,II22771,II22802
	,II22833,II22864,II22895,II22926,II22957,II22988,II26020,II26051
	,II26082,II26113,II26144,II26175,II26206,II26237,II26268,II26299
	,II26330,II26361,II26392,II26423,II26454,II26485,II26516,II26547
	,II26578,II26609,II26640,II26671,II26702,II26733,II26764,II26795
	,II26826,II26857,II26888,II26919,II26950,II26981,II26032,II26063
	,II26094,II26125,II26156,II26187,II26218,II26249,II26280,II26311
	,II26342,II26373,II26404,II26435,II26466,II26497,II26528,II26559
	,II26590,II26621,II26652,II26683,II26714,II26745,II26776,II26807
	,II26838,II26869,II26900,II26931,II26962,II26993,II30025,II30056
	,II30087,II30118,II30149,II30180,II30211,II30242,II30273,II30304
	,II30335,II30366,II30397,II30428,II30459,II30490,II30521,II30552
	,II30583,II30614,II30645,II30676,II30707,II30738,II30769,II30800
	,II30831,II30862,II30893,II30924,II30955,II30986,II30037,II30068
	,II30099,II30130,II30161,II30192,II30223,II30254,II30285,II30316
	,II30347,II30378,II30409,II30440,II30471,II30502,II30533,II30564
	,II30595,II30626,II30657,II30688,II30719,II30750,II30781,II30812
	,II30843,II30874,II30905,II30936,II30967,II30998,II34030,II34061
	,II34092,II34123,II34154,II34185,II34216,II34247,II34278,II34309
	,II34340,II34371,II34402,II34433,II34464,II34495,II34526,II34557
	,II34588,II34619,II34650,II34681,II34712,II34743,II34774,II34805
	,II34836,II34867,II34898,II34929,II34960,II34991,II34042,II34073
	,II34104,II34135,II34166,II34197,II34228,II34259,II34290,II34321
	,II34352,II34383,II34414,II34445,II34476,II34507,II34538,II34569
	,II34600,II34631,II34662,II34693,II34724,II34755,II34786,II34817
	,II34848,II34879,II34910,II34941,II34972,II35003,II35555,II35751
	,II35744,II35737,II35541,II35730,II35723,II35716,II35709,II35702
	,II35695,II35526,II35688,II35681,II35674,II35667,II35511,II35660
	,II35653,II35646,II35639,II35632,II35625,II35618,II35611,II35604
	,II35597,II35590,II35583,II35576,II35569,II35562,II31550,II31746
	,II31739,II31732,II31536,II31725,II31718,II31711,II31704,II31697
	,II31690,II31521,II31683,II31676,II31669,II31662,II31506,II31655
	,II31648,II31641,II31634,II31627,II31620,II31613,II31606,II31599
	,II31592,II31585,II31578,II31571,II31564,II31557,II27545,II27741
	,II27734,II27727,II27531,II27720,II27713,II27706,II27699,II27692
	,II27685,II27516,II27678,II27671,II27664,II27657,II27501,II27650
	,II27643,II27636,II27629,II27622,II27615,II27608,II27601,II27594
	,II27587,II27580,II27573,II27566,II27559,II27552,II23540,II23736
	,II23729,II23722,II23526,II23715,II23708,II23701,II23694,II23687
	,II23680,II23511,II23673,II23666,II23659,II23652,II23496,II23645
	,II23638,II23631,II23624,II23617,II23610,II23603,II23596,II23589
	,II23582,II23575,II23568,II23561,II23554,II23547,II19535,II19731
	,II19724,II19717,II19521,II19710,II19703,II19696,II19689,II19682
	,II19675,II19506,II19668,II19661,II19654,II19647,II19491,II19640
	,II19633,II19626,II19619,II19612,II19605,II19598,II19591,II19584
	,II19577,II19570,II19563,II19556,II19549,II19542,II15530,II15726
	,II15719,II15712,II15516,II15705,II15698,II15691,II15684,II15677
	,II15670,II15501,II15663,II15656,II15649,II15642,II15486,II15635
	,II15628,II15621,II15614,II15607,II15600,II15593,II15586,II15579
	,II15572,II15565,II15558,II15551,II15544,II15537,II11525,II11721
	,II11714,II11707,II11511,II11700,II11693,II11686,II11679,II11672
	,II11665,II11496,II11658,II11651,II11644,II11637,II11481,II11630
	,II11623,II11616,II11609,II11602,II11595,II11588,II11581,II11574
	,II11567,II11560,II11553,II11546,II11539,II11532,II7520,II7716
	,II7709,II7702,II7506,II7695,II7688,II7681,II7674,II7667
	,II7660,II7491,II7653,II7646,II7639,II7632,II7476,II7625
	,II7618,II7611,II7604,II7597,II7590,II7583,II7576,II7569
	,II7562,II7555,II7548,II7541,II7534,II7527,II3515,II3711
	,II3704,II3697,II3501,II3690,II3683,II3676,II3669,II3662
	,II3655,II3486,II3648,II3641,II3634,II3627,II3471,II3620
	,II3613,II3606,II3599,II3592,II3585,II3578,II3571,II3564
	,II3557,II3550,II3543,II3536,II3529,II3522,II3712,II3705
	,II3698,II3691,II3684,II3677,II3670,II3663,II3656,II3649
	,II3642,II3635,II3628,II3621,II3614,II3607,II3600,II3593
	,II3586,II3579,II3572,II3565,II3558,II3551,II3544,II3537
	,II3530,II3523,II3516,II3502,II3487,II3472,II7717,II7710
	,II7703,II7696,II7689,II7682,II7675,II7668,II7661,II7654
	,II7647,II7640,II7633,II7626,II7619,II7612,II7605,II7598
	,II7591,II7584,II7577,II7570,II7563,II7556,II7549,II7542
	,II7535,II7528,II7521,II7507,II7492,II7477,II11722,II11715
	,II11708,II11701,II11694,II11687,II11680,II11673,II11666,II11659
	,II11652,II11645,II11638,II11631,II11624,II11617,II11610,II11603
	,II11596,II11589,II11582,II11575,II11568,II11561,II11554,II11547
	,II11540,II11533,II11526,II11512,II11497,II11482,II15727,II15720
	,II15713,II15706,II15699,II15692,II15685,II15678,II15671,II15664
	,II15657,II15650,II15643,II15636,II15629,II15622,II15615,II15608
	,II15601,II15594,II15587,II15580,II15573,II15566,II15559,II15552
	,II15545,II15538,II15531,II15517,II15502,II15487,II19732,II19725
	,II19718,II19711,II19704,II19697,II19690,II19683,II19676,II19669
	,II19662,II19655,II19648,II19641,II19634,II19627,II19620,II19613
	,II19606,II19599,II19592,II19585,II19578,II19571,II19564,II19557
	,II19550,II19543,II19536,II19522,II19507,II19492,II23737,II23730
	,II23723,II23716,II23709,II23702,II23695,II23688,II23681,II23674
	,II23667,II23660,II23653,II23646,II23639,II23632,II23625,II23618
	,II23611,II23604,II23597,II23590,II23583,II23576,II23569,II23562
	,II23555,II23548,II23541,II23527,II23512,II23497,II27742,II27735
	,II27728,II27721,II27714,II27707,II27700,II27693,II27686,II27679
	,II27672,II27665,II27658,II27651,II27644,II27637,II27630,II27623
	,II27616,II27609,II27602,II27595,II27588,II27581,II27574,II27567
	,II27560,II27553,II27546,II27532,II27517,II27502,II31747,II31740
	,II31733,II31726,II31719,II31712,II31705,II31698,II31691,II31684
	,II31677,II31670,II31663,II31656,II31649,II31642,II31635,II31628
	,II31621,II31614,II31607,II31600,II31593,II31586,II31579,II31572
	,II31565,II31558,II31551,II31537,II31522,II31507,II35752,II35745
	,II35738,II35731,II35724,II35717,II35710,II35703,II35696,II35689
	,II35682,II35675,II35668,II35661,II35654,II35647,II35640,II35633
	,II35626,II35619,II35612,II35605,II35598,II35591,II35584,II35577
	,II35570,II35563,II35556,II35542,II35527,II35512,II34988,II34957
	,II34926,II34895,II34864,II34833,II34802,II34771,II34740,II34709
	,II34678,II34647,II34616,II34585,II34554,II34523,II34492,II34461
	,II34430,II34399,II34368,II34337,II34306,II34275,II34244,II34213
	,II34182,II34151,II34120,II34089,II34058,II34027,II30983,II30952
	,II30921,II30890,II30859,II30828,II30797,II30766,II30735,II30704
	,II30673,II30642,II30611,II30580,II30549,II30518,II30487,II30456
	,II30425,II30394,II30363,II30332,II30301,II30270,II30239,II30208
	,II30177,II30146,II30115,II30084,II30053,II30022,II26978,II26947
	,II26916,II26885,II26854,II26823,II26792,II26761,II26730,II26699
	,II26668,II26637,II26606,II26575,II26544,II26513,II26482,II26451
	,II26420,II26389,II26358,II26327,II26296,II26265,II26234,II26203
	,II26172,II26141,II26110,II26079,II26048,II26017,II22973,II22942
	,II22911,II22880,II22849,II22818,II22787,II22756,II22725,II22694
	,II22663,II22632,II22601,II22570,II22539,II22508,II22477,II22446
	,II22415,II22384,II22353,II22322,II22291,II22260,II22229,II22198
	,II22167,II22136,II22105,II22074,II22043,II22012,II18968,II18937
	,II18906,II18875,II18844,II18813,II18782,II18751,II18720,II18689
	,II18658,II18627,II18596,II18565,II18534,II18503,II18472,II18441
	,II18410,II18379,II18348,II18317,II18286,II18255,II18224,II18193
	,II18162,II18131,II18100,II18069,II18038,II18007,II14963,II14932
	,II14901,II14870,II14839,II14808,II14777,II14746,II14715,II14684
	,II14653,II14622,II14591,II14560,II14529,II14498,II14467,II14436
	,II14405,II14374,II14343,II14312,II14281,II14250,II14219,II14188
	,II14157,II14126,II14095,II14064,II14033,II14002,II10958,II10927
	,II10896,II10865,II10834,II10803,II10772,II10741,II10710,II10679
	,II10648,II10617,II10586,II10555,II10524,II10493,II10462,II10431
	,II10400,II10369,II10338,II10307,II10276,II10245,II10214,II10183
	,II10152,II10121,II10090,II10059,II10028,II9997,II6953,II6922
	,II6891,II6860,II6829,II6798,II6767,II6736,II6705,II6674
	,II6643,II6612,II6581,II6550,II6519,II6488,II6457,II6426
	,II6395,II6364,II6333,II6302,II6271,II6240,II6209,II6178
	,II6147,II6116,II6085,II6054,II6023,II5992,II2948,II2917
	,II2886,II2855,II2824,II2793,II2762,II2731,II2700,II2669
	,II2638,II2607,II2576,II2545,II2514,II2483,II2452,II2421
	,II2390,II2359,II2328,II2297,II2266,II2235,II2204,II2173
	,II2142,II2111,II2080,II2049,II2018,II1987,WX10386,WX10400
	,WX10414,WX10428,WX10442,WX10456,WX10470,WX10484,WX10498,WX10512
	,WX10526,WX10540,WX10554,WX10568,WX10582,WX10596,WX10610,WX10624
	,WX10638,WX10652,WX10666,WX10680,WX10694,WX10708,WX10722,WX10736
	,WX10750,WX10764,WX10778,WX10792,WX10806,WX10820,WX1262,WX1261
	,WX1260,WX1259,WX1258,WX1257,WX1256,WX1255,WX1254,WX1253
	,WX1252,WX1251,WX1250,WX1249,WX1248,WX1247,WX1246,WX1245
	,WX1244,WX1243,WX1242,WX1241,WX1240,WX1239,WX1238,WX1237
	,WX1236,WX1235,WX1234,II3499,II3484,II3469,WX2555,WX2554
	,WX2553,WX2552,WX2551,WX2550,WX2549,WX2548,WX2547,WX2546
	,WX2545,WX2544,WX2543,WX2542,WX2541,WX2540,WX2539,WX2538
	,WX2537,WX2536,WX2535,WX2534,WX2533,WX2532,WX2531,WX2530
	,WX2529,WX2528,WX2527,II7504,II7489,II7474,WX3848,WX3847
	,WX3846,WX3845,WX3844,WX3843,WX3842,WX3841,WX3840,WX3839
	,WX3838,WX3837,WX3836,WX3835,WX3834,WX3833,WX3832,WX3831
	,WX3830,WX3829,WX3828,WX3827,WX3826,WX3825,WX3824,WX3823
	,WX3822,WX3821,WX3820,II11509,II11494,II11479,WX5141,WX5140
	,WX5139,WX5138,WX5137,WX5136,WX5135,WX5134,WX5133,WX5132
	,WX5131,WX5130,WX5129,WX5128,WX5127,WX5126,WX5125,WX5124
	,WX5123,WX5122,WX5121,WX5120,WX5119,WX5118,WX5117,WX5116
	,WX5115,WX5114,WX5113,II15514,II15499,II15484,WX6434,WX6433
	,WX6432,WX6431,WX6430,WX6429,WX6428,WX6427,WX6426,WX6425
	,WX6424,WX6423,WX6422,WX6421,WX6420,WX6419,WX6418,WX6417
	,WX6416,WX6415,WX6414,WX6413,WX6412,WX6411,WX6410,WX6409
	,WX6408,WX6407,WX6406,II19519,II19504,II19489,WX7727,WX7726
	,WX7725,WX7724,WX7723,WX7722,WX7721,WX7720,WX7719,WX7718
	,WX7717,WX7716,WX7715,WX7714,WX7713,WX7712,WX7711,WX7710
	,WX7709,WX7708,WX7707,WX7706,WX7705,WX7704,WX7703,WX7702
	,WX7701,WX7700,WX7699,II23524,II23509,II23494,WX9020,WX9019
	,WX9018,WX9017,WX9016,WX9015,WX9014,WX9013,WX9012,WX9011
	,WX9010,WX9009,WX9008,WX9007,WX9006,WX9005,WX9004,WX9003
	,WX9002,WX9001,WX9000,WX8999,WX8998,WX8997,WX8996,WX8995
	,WX8994,WX8993,WX8992,II27529,II27514,II27499,WX10313,WX10312
	,WX10311,WX10310,WX10309,WX10308,WX10307,WX10306,WX10305,WX10304
	,WX10303,WX10302,WX10301,WX10300,WX10299,WX10298,WX10297,WX10296
	,WX10295,WX10294,WX10293,WX10292,WX10291,WX10290,WX10289,WX10288
	,WX10287,WX10286,WX10285,II31534,II31519,II31504,WX11606,WX11605
	,WX11604,WX11603,WX11602,WX11601,WX11600,WX11599,WX11598,WX11597
	,WX11596,WX11595,WX11594,WX11593,WX11592,WX11591,WX11590,WX11589
	,WX11588,WX11587,WX11586,WX11585,WX11584,WX11583,WX11582,WX11581
	,WX11580,WX11579,WX11578,II35539,II35524,II35509,WX10814,WX10800
	,WX10786,WX10772,WX10758,WX10744,WX10730,WX10716,WX10702,WX10688
	,WX10674,WX10660,WX10646,WX10632,WX10618,WX10604,WX10590,WX10576
	,WX10562,WX10548,WX10534,WX10520,WX10506,WX10492,WX10478,WX10464
	,WX10450,WX10436,WX10422,WX10408,WX10394,WX10380,II34996,II34965
	,II34934,II34903,II34872,II34841,II34810,II34779,II34748,II34717
	,II34686,II34655,II34624,II34593,II34562,II34531,II34500,II34469
	,II34438,II34407,II34376,II34345,II34314,II34283,II34252,II34221
	,II34190,II34159,II34128,II34097,II34066,II34035,II30991,II30960
	,II30929,II30898,II30867,II30836,II30805,II30774,II30743,II30712
	,II30681,II30650,II30619,II30588,II30557,II30526,II30495,II30464
	,II30433,II30402,II30371,II30340,II30309,II30278,II30247,II30216
	,II30185,II30154,II30123,II30092,II30061,II30030,II26986,II26955
	,II26924,II26893,II26862,II26831,II26800,II26769,II26738,II26707
	,II26676,II26645,II26614,II26583,II26552,II26521,II26490,II26459
	,II26428,II26397,II26366,II26335,II26304,II26273,II26242,II26211
	,II26180,II26149,II26118,II26087,II26056,II26025,II22981,II22950
	,II22919,II22888,II22857,II22826,II22795,II22764,II22733,II22702
	,II22671,II22640,II22609,II22578,II22547,II22516,II22485,II22454
	,II22423,II22392,II22361,II22330,II22299,II22268,II22237,II22206
	,II22175,II22144,II22113,II22082,II22051,II22020,II18976,II18945
	,II18914,II18883,II18852,II18821,II18790,II18759,II18728,II18697
	,II18666,II18635,II18604,II18573,II18542,II18511,II18480,II18449
	,II18418,II18387,II18356,II18325,II18294,II18263,II18232,II18201
	,II18170,II18139,II18108,II18077,II18046,II18015,II14971,II14940
	,II14909,II14878,II14847,II14816,II14785,II14754,II14723,II14692
	,II14661,II14630,II14599,II14568,II14537,II14506,II14475,II14444
	,II14413,II14382,II14351,II14320,II14289,II14258,II14227,II14196
	,II14165,II14134,II14103,II14072,II14041,II14010,II10966,II10935
	,II10904,II10873,II10842,II10811,II10780,II10749,II10718,II10687
	,II10656,II10625,II10594,II10563,II10532,II10501,II10470,II10439
	,II10408,II10377,II10346,II10315,II10284,II10253,II10222,II10191
	,II10160,II10129,II10098,II10067,II10036,II10005,II6961,II6930
	,II6899,II6868,II6837,II6806,II6775,II6744,II6713,II6682
	,II6651,II6620,II6589,II6558,II6527,II6496,II6465,II6434
	,II6403,II6372,II6341,II6310,II6279,II6248,II6217,II6186
	,II6155,II6124,II6093,II6062,II6031,II6000,II2956,II2925
	,II2894,II2863,II2832,II2801,II2770,II2739,II2708,II2677
	,II2646,II2615,II2584,II2553,II2522,II2491,II2460,II2429
	,II2398,II2367,II2336,II2305,II2274,II2243,II2212,II2181
	,II2150,II2119,II2088,II2057,II2026,II1995,WX11670,WX11668
	,WX11666,WX11664,WX11662,WX11660,WX11658,WX11656,WX11654,WX11652
	,WX11650,WX11648,WX11646,WX11644,WX11642,WX11638,WX11636,WX11634
	,WX11632,WX11628,WX11626,WX11624,WX11622,WX11620,WX11618,WX11614
	,WX11612,WX11610,WX11608,WX10377,WX10375,WX10373,WX10371,WX10369
	,WX10367,WX10365,WX10363,WX10361,WX10359,WX10357,WX10355,WX10353
	,WX10351,WX10349,WX10345,WX10343,WX10341,WX10339,WX10335,WX10333
	,WX10331,WX10329,WX10327,WX10325,WX10321,WX10319,WX10317,WX10315
	,WX9084,WX9082,WX9080,WX9078,WX9076,WX9074,WX9072,WX9070
	,WX9068,WX9066,WX9064,WX9062,WX9060,WX9058,WX9056,WX9052
	,WX9050,WX9048,WX9046,WX9042,WX9040,WX9038,WX9036,WX9034
	,WX9032,WX9028,WX9026,WX9024,WX9022,WX7791,WX7789,WX7787
	,WX7785,WX7783,WX7781,WX7779,WX7777,WX7775,WX7773,WX7771
	,WX7769,WX7767,WX7765,WX7763,WX7759,WX7757,WX7755,WX7753
	,WX7749,WX7747,WX7745,WX7743,WX7741,WX7739,WX7735,WX7733
	,WX7731,WX7729,WX6498,WX6496,WX6494,WX6492,WX6490,WX6488
	,WX6486,WX6484,WX6482,WX6480,WX6478,WX6476,WX6474,WX6472
	,WX6470,WX6466,WX6464,WX6462,WX6460,WX6456,WX6454,WX6452
	,WX6450,WX6448,WX6446,WX6442,WX6440,WX6438,WX6436,WX5205
	,WX5203,WX5201,WX5199,WX5197,WX5195,WX5193,WX5191,WX5189
	,WX5187,WX5185,WX5183,WX5181,WX5179,WX5177,WX5173,WX5171
	,WX5169,WX5167,WX5163,WX5161,WX5159,WX5157,WX5155,WX5153
	,WX5149,WX5147,WX5145,WX5143,WX3912,WX3910,WX3908,WX3906
	,WX3904,WX3902,WX3900,WX3898,WX3896,WX3894,WX3892,WX3890
	,WX3888,WX3886,WX3884,WX3880,WX3878,WX3876,WX3874,WX3870
	,WX3868,WX3866,WX3864,WX3862,WX3860,WX3856,WX3854,WX3852
	,WX3850,WX2619,WX2617,WX2615,WX2613,WX2611,WX2609,WX2607
	,WX2605,WX2603,WX2601,WX2599,WX2597,WX2595,WX2593,WX2591
	,WX2587,WX2585,WX2583,WX2581,WX2577,WX2575,WX2573,WX2571
	,WX2569,WX2567,WX2563,WX2561,WX2559,WX2557,WX1326,WX1324
	,WX1322,WX1320,WX1318,WX1316,WX1314,WX1312,WX1310,WX1308
	,WX1306,WX1304,WX1302,WX1300,WX1298,WX1294,WX1292,WX1290
	,WX1288,WX1284,WX1282,WX1280,WX1278,WX1276,WX1274,WX1270
	,WX1268,WX1266,WX1264,II3507,II3492,II3477,II7512,II7497
	,II7482,II11517,II11502,II11487,II15522,II15507,II15492,II19527
	,II19512,II19497,II23532,II23517,II23502,II27537,II27522,II27507
	,II31542,II31527,II31512,II35547,II35532,II35517,II1997,II2028
	,II2059,II2090,II2121,II2152,II2183,II2214,II2245,II2276
	,II2307,II2338,II2369,II2400,II2431,II2462,II2493,II2524
	,II2555,II2586,II2617,II2648,II2679,II2710,II2741,II2772
	,II2803,II2834,II2865,II2896,II2927,II2958,II1996,II2027
	,II2058,II2089,II2120,II2151,II2182,II2213,II2244,II2275
	,II2306,II2337,II2368,II2399,II2430,II2461,II2492,II2523
	,II2554,II2585,II2616,II2647,II2678,II2709,II2740,II2771
	,II2802,II2833,II2864,II2895,II2926,II2957,II6002,II6033
	,II6064,II6095,II6126,II6157,II6188,II6219,II6250,II6281
	,II6312,II6343,II6374,II6405,II6436,II6467,II6498,II6529
	,II6560,II6591,II6622,II6653,II6684,II6715,II6746,II6777
	,II6808,II6839,II6870,II6901,II6932,II6963,II6001,II6032
	,II6063,II6094,II6125,II6156,II6187,II6218,II6249,II6280
	,II6311,II6342,II6373,II6404,II6435,II6466,II6497,II6528
	,II6559,II6590,II6621,II6652,II6683,II6714,II6745,II6776
	,II6807,II6838,II6869,II6900,II6931,II6962,II10007,II10038
	,II10069,II10100,II10131,II10162,II10193,II10224,II10255,II10286
	,II10317,II10348,II10379,II10410,II10441,II10472,II10503,II10534
	,II10565,II10596,II10627,II10658,II10689,II10720,II10751,II10782
	,II10813,II10844,II10875,II10906,II10937,II10968,II10006,II10037
	,II10068,II10099,II10130,II10161,II10192,II10223,II10254,II10285
	,II10316,II10347,II10378,II10409,II10440,II10471,II10502,II10533
	,II10564,II10595,II10626,II10657,II10688,II10719,II10750,II10781
	,II10812,II10843,II10874,II10905,II10936,II10967,II14012,II14043
	,II14074,II14105,II14136,II14167,II14198,II14229,II14260,II14291
	,II14322,II14353,II14384,II14415,II14446,II14477,II14508,II14539
	,II14570,II14601,II14632,II14663,II14694,II14725,II14756,II14787
	,II14818,II14849,II14880,II14911,II14942,II14973,II14011,II14042
	,II14073,II14104,II14135,II14166,II14197,II14228,II14259,II14290
	,II14321,II14352,II14383,II14414,II14445,II14476,II14507,II14538
	,II14569,II14600,II14631,II14662,II14693,II14724,II14755,II14786
	,II14817,II14848,II14879,II14910,II14941,II14972,II18017,II18048
	,II18079,II18110,II18141,II18172,II18203,II18234,II18265,II18296
	,II18327,II18358,II18389,II18420,II18451,II18482,II18513,II18544
	,II18575,II18606,II18637,II18668,II18699,II18730,II18761,II18792
	,II18823,II18854,II18885,II18916,II18947,II18978,II18016,II18047
	,II18078,II18109,II18140,II18171,II18202,II18233,II18264,II18295
	,II18326,II18357,II18388,II18419,II18450,II18481,II18512,II18543
	,II18574,II18605,II18636,II18667,II18698,II18729,II18760,II18791
	,II18822,II18853,II18884,II18915,II18946,II18977,II22022,II22053
	,II22084,II22115,II22146,II22177,II22208,II22239,II22270,II22301
	,II22332,II22363,II22394,II22425,II22456,II22487,II22518,II22549
	,II22580,II22611,II22642,II22673,II22704,II22735,II22766,II22797
	,II22828,II22859,II22890,II22921,II22952,II22983,II22021,II22052
	,II22083,II22114,II22145,II22176,II22207,II22238,II22269,II22300
	,II22331,II22362,II22393,II22424,II22455,II22486,II22517,II22548
	,II22579,II22610,II22641,II22672,II22703,II22734,II22765,II22796
	,II22827,II22858,II22889,II22920,II22951,II22982,II26027,II26058
	,II26089,II26120,II26151,II26182,II26213,II26244,II26275,II26306
	,II26337,II26368,II26399,II26430,II26461,II26492,II26523,II26554
	,II26585,II26616,II26647,II26678,II26709,II26740,II26771,II26802
	,II26833,II26864,II26895,II26926,II26957,II26988,II26026,II26057
	,II26088,II26119,II26150,II26181,II26212,II26243,II26274,II26305
	,II26336,II26367,II26398,II26429,II26460,II26491,II26522,II26553
	,II26584,II26615,II26646,II26677,II26708,II26739,II26770,II26801
	,II26832,II26863,II26894,II26925,II26956,II26987,II30032,II30063
	,II30094,II30125,II30156,II30187,II30218,II30249,II30280,II30311
	,II30342,II30373,II30404,II30435,II30466,II30497,II30528,II30559
	,II30590,II30621,II30652,II30683,II30714,II30745,II30776,II30807
	,II30838,II30869,II30900,II30931,II30962,II30993,II30031,II30062
	,II30093,II30124,II30155,II30186,II30217,II30248,II30279,II30310
	,II30341,II30372,II30403,II30434,II30465,II30496,II30527,II30558
	,II30589,II30620,II30651,II30682,II30713,II30744,II30775,II30806
	,II30837,II30868,II30899,II30930,II30961,II30992,II34037,II34068
	,II34099,II34130,II34161,II34192,II34223,II34254,II34285,II34316
	,II34347,II34378,II34409,II34440,II34471,II34502,II34533,II34564
	,II34595,II34626,II34657,II34688,II34719,II34750,II34781,II34812
	,II34843,II34874,II34905,II34936,II34967,II34998,II34036,II34067
	,II34098,II34129,II34160,II34191,II34222,II34253,II34284,II34315
	,II34346,II34377,II34408,II34439,II34470,II34501,II34532,II34563
	,II34594,II34625,II34656,II34687,II34718,II34749,II34780,II34811
	,II34842,II34873,II34904,II34935,II34966,II34997,II35519,II35534
	,II35549,II31514,II31529,II31544,II27509,II27524,II27539,II23504
	,II23519,II23534,II19499,II19514,II19529,II15494,II15509,II15524
	,II11489,II11504,II11519,II7484,II7499,II7514,II3479,II3494
	,II3509,II3508,II3493,II3478,II7513,II7498,II7483,II11518
	,II11503,II11488,II15523,II15508,II15493,II19528,II19513,II19498
	,II23533,II23518,II23503,II27538,II27523,II27508,II31543,II31528
	,II31513,II35548,II35533,II35518,II34987,II34956,II34925,II34894
	,II34863,II34832,II34801,II34770,II34739,II34708,II34677,II34646
	,II34615,II34584,II34553,II34522,II34491,II34460,II34429,II34398
	,II34367,II34336,II34305,II34274,II34243,II34212,II34181,II34150
	,II34119,II34088,II34057,II34026,II30982,II30951,II30920,II30889
	,II30858,II30827,II30796,II30765,II30734,II30703,II30672,II30641
	,II30610,II30579,II30548,II30517,II30486,II30455,II30424,II30393
	,II30362,II30331,II30300,II30269,II30238,II30207,II30176,II30145
	,II30114,II30083,II30052,II30021,II26977,II26946,II26915,II26884
	,II26853,II26822,II26791,II26760,II26729,II26698,II26667,II26636
	,II26605,II26574,II26543,II26512,II26481,II26450,II26419,II26388
	,II26357,II26326,II26295,II26264,II26233,II26202,II26171,II26140
	,II26109,II26078,II26047,II26016,II22972,II22941,II22910,II22879
	,II22848,II22817,II22786,II22755,II22724,II22693,II22662,II22631
	,II22600,II22569,II22538,II22507,II22476,II22445,II22414,II22383
	,II22352,II22321,II22290,II22259,II22228,II22197,II22166,II22135
	,II22104,II22073,II22042,II22011,II18967,II18936,II18905,II18874
	,II18843,II18812,II18781,II18750,II18719,II18688,II18657,II18626
	,II18595,II18564,II18533,II18502,II18471,II18440,II18409,II18378
	,II18347,II18316,II18285,II18254,II18223,II18192,II18161,II18130
	,II18099,II18068,II18037,II18006,II14962,II14931,II14900,II14869
	,II14838,II14807,II14776,II14745,II14714,II14683,II14652,II14621
	,II14590,II14559,II14528,II14497,II14466,II14435,II14404,II14373
	,II14342,II14311,II14280,II14249,II14218,II14187,II14156,II14125
	,II14094,II14063,II14032,II14001,II10957,II10926,II10895,II10864
	,II10833,II10802,II10771,II10740,II10709,II10678,II10647,II10616
	,II10585,II10554,II10523,II10492,II10461,II10430,II10399,II10368
	,II10337,II10306,II10275,II10244,II10213,II10182,II10151,II10120
	,II10089,II10058,II10027,II9996,II6952,II6921,II6890,II6859
	,II6828,II6797,II6766,II6735,II6704,II6673,II6642,II6611
	,II6580,II6549,II6518,II6487,II6456,II6425,II6394,II6363
	,II6332,II6301,II6270,II6239,II6208,II6177,II6146,II6115
	,II6084,II6053,II6022,II5991,II2947,II2916,II2885,II2854
	,II2823,II2792,II2761,II2730,II2699,II2668,II2637,II2606
	,II2575,II2544,II2513,II2482,II2451,II2420,II2389,II2358
	,II2327,II2296,II2265,II2234,II2203,II2172,II2141,II2110
	,II2079,II2048,II2017,II1986,WX1233,WX1232,WX1231,WX2526
	,WX2525,WX2524,WX3819,WX3818,WX3817,WX5112,WX5111,WX5110
	,WX6405,WX6404,WX6403,WX7698,WX7697,WX7696,WX8991,WX8990
	,WX8989,WX10284,WX10283,WX10282,WX11577,WX11576,WX11575,II35011
	,II34980,II34949,II34918,II34887,II34856,II34825,II34794,II34763
	,II34732,II34701,II34670,II34639,II34608,II34577,II34546,II34515
	,II34484,II34453,II34422,II34391,II34360,II34329,II34298,II34267
	,II34236,II34205,II34174,II34143,II34112,II34081,II34050,II31006
	,II30975,II30944,II30913,II30882,II30851,II30820,II30789,II30758
	,II30727,II30696,II30665,II30634,II30603,II30572,II30541,II30510
	,II30479,II30448,II30417,II30386,II30355,II30324,II30293,II30262
	,II30231,II30200,II30169,II30138,II30107,II30076,II30045,II27001
	,II26970,II26939,II26908,II26877,II26846,II26815,II26784,II26753
	,II26722,II26691,II26660,II26629,II26598,II26567,II26536,II26505
	,II26474,II26443,II26412,II26381,II26350,II26319,II26288,II26257
	,II26226,II26195,II26164,II26133,II26102,II26071,II26040,II22996
	,II22965,II22934,II22903,II22872,II22841,II22810,II22779,II22748
	,II22717,II22686,II22655,II22624,II22593,II22562,II22531,II22500
	,II22469,II22438,II22407,II22376,II22345,II22314,II22283,II22252
	,II22221,II22190,II22159,II22128,II22097,II22066,II22035,II18991
	,II18960,II18929,II18898,II18867,II18836,II18805,II18774,II18743
	,II18712,II18681,II18650,II18619,II18588,II18557,II18526,II18495
	,II18464,II18433,II18402,II18371,II18340,II18309,II18278,II18247
	,II18216,II18185,II18154,II18123,II18092,II18061,II18030,II14986
	,II14955,II14924,II14893,II14862,II14831,II14800,II14769,II14738
	,II14707,II14676,II14645,II14614,II14583,II14552,II14521,II14490
	,II14459,II14428,II14397,II14366,II14335,II14304,II14273,II14242
	,II14211,II14180,II14149,II14118,II14087,II14056,II14025,II10981
	,II10950,II10919,II10888,II10857,II10826,II10795,II10764,II10733
	,II10702,II10671,II10640,II10609,II10578,II10547,II10516,II10485
	,II10454,II10423,II10392,II10361,II10330,II10299,II10268,II10237
	,II10206,II10175,II10144,II10113,II10082,II10051,II10020,II6976
	,II6945,II6914,II6883,II6852,II6821,II6790,II6759,II6728
	,II6697,II6666,II6635,II6604,II6573,II6542,II6511,II6480
	,II6449,II6418,II6387,II6356,II6325,II6294,II6263,II6232
	,II6201,II6170,II6139,II6108,II6077,II6046,II6015,II2971
	,II2940,II2909,II2878,II2847,II2816,II2785,II2754,II2723
	,II2692,II2661,II2630,II2599,II2568,II2537,II2506,II2475
	,II2444,II2413,II2382,II2351,II2320,II2289,II2258,II2227
	,II2196,II2165,II2134,II2103,II2072,II2041,II2010,WX11640
	,WX11630,WX11616,WX10347,WX10337,WX10323,WX9054,WX9044,WX9030
	,WX7761,WX7751,WX7737,WX6468,WX6458,WX6444,WX5175,WX5165
	,WX5151,WX3882,WX3872,WX3858,WX2589,WX2579,WX2565,WX1296
	,WX1286,WX1272,II2011,II2042,II2073,II2104,II2135,II2166
	,II2197,II2228,II2259,II2290,II2321,II2352,II2383,II2414
	,II2445,II2476,II2507,II2538,II2569,II2600,II2631,II2662
	,II2693,II2724,II2755,II2786,II2817,II2848,II2879,II2910
	,II2941,II2972,II6016,II6047,II6078,II6109,II6140,II6171
	,II6202,II6233,II6264,II6295,II6326,II6357,II6388,II6419
	,II6450,II6481,II6512,II6543,II6574,II6605,II6636,II6667
	,II6698,II6729,II6760,II6791,II6822,II6853,II6884,II6915
	,II6946,II6977,II10021,II10052,II10083,II10114,II10145,II10176
	,II10207,II10238,II10269,II10300,II10331,II10362,II10393,II10424
	,II10455,II10486,II10517,II10548,II10579,II10610,II10641,II10672
	,II10703,II10734,II10765,II10796,II10827,II10858,II10889,II10920
	,II10951,II10982,II14026,II14057,II14088,II14119,II14150,II14181
	,II14212,II14243,II14274,II14305,II14336,II14367,II14398,II14429
	,II14460,II14491,II14522,II14553,II14584,II14615,II14646,II14677
	,II14708,II14739,II14770,II14801,II14832,II14863,II14894,II14925
	,II14956,II14987,II18031,II18062,II18093,II18124,II18155,II18186
	,II18217,II18248,II18279,II18310,II18341,II18372,II18403,II18434
	,II18465,II18496,II18527,II18558,II18589,II18620,II18651,II18682
	,II18713,II18744,II18775,II18806,II18837,II18868,II18899,II18930
	,II18961,II18992,II22036,II22067,II22098,II22129,II22160,II22191
	,II22222,II22253,II22284,II22315,II22346,II22377,II22408,II22439
	,II22470,II22501,II22532,II22563,II22594,II22625,II22656,II22687
	,II22718,II22749,II22780,II22811,II22842,II22873,II22904,II22935
	,II22966,II22997,II26041,II26072,II26103,II26134,II26165,II26196
	,II26227,II26258,II26289,II26320,II26351,II26382,II26413,II26444
	,II26475,II26506,II26537,II26568,II26599,II26630,II26661,II26692
	,II26723,II26754,II26785,II26816,II26847,II26878,II26909,II26940
	,II26971,II27002,II30046,II30077,II30108,II30139,II30170,II30201
	,II30232,II30263,II30294,II30325,II30356,II30387,II30418,II30449
	,II30480,II30511,II30542,II30573,II30604,II30635,II30666,II30697
	,II30728,II30759,II30790,II30821,II30852,II30883,II30914,II30945
	,II30976,II31007,II34051,II34082,II34113,II34144,II34175,II34206
	,II34237,II34268,II34299,II34330,II34361,II34392,II34423,II34454
	,II34485,II34516,II34547,II34578,II34609,II34640,II34671,II34702
	,II34733,II34764,II34795,II34826,II34857,II34888,II34919,II34950
	,II34981,II35012,II35013,II34982,II34951,II34920,II34889,II34858
	,II34827,II34796,II34765,II34734,II34703,II34672,II34641,II34610
	,II34579,II34548,II34517,II34486,II34455,II34424,II34393,II34362
	,II34331,II34300,II34269,II34238,II34207,II34176,II34145,II34114
	,II34083,II34052,II31008,II30977,II30946,II30915,II30884,II30853
	,II30822,II30791,II30760,II30729,II30698,II30667,II30636,II30605
	,II30574,II30543,II30512,II30481,II30450,II30419,II30388,II30357
	,II30326,II30295,II30264,II30233,II30202,II30171,II30140,II30109
	,II30078,II30047,II27003,II26972,II26941,II26910,II26879,II26848
	,II26817,II26786,II26755,II26724,II26693,II26662,II26631,II26600
	,II26569,II26538,II26507,II26476,II26445,II26414,II26383,II26352
	,II26321,II26290,II26259,II26228,II26197,II26166,II26135,II26104
	,II26073,II26042,II22998,II22967,II22936,II22905,II22874,II22843
	,II22812,II22781,II22750,II22719,II22688,II22657,II22626,II22595
	,II22564,II22533,II22502,II22471,II22440,II22409,II22378,II22347
	,II22316,II22285,II22254,II22223,II22192,II22161,II22130,II22099
	,II22068,II22037,II18993,II18962,II18931,II18900,II18869,II18838
	,II18807,II18776,II18745,II18714,II18683,II18652,II18621,II18590
	,II18559,II18528,II18497,II18466,II18435,II18404,II18373,II18342
	,II18311,II18280,II18249,II18218,II18187,II18156,II18125,II18094
	,II18063,II18032,II14988,II14957,II14926,II14895,II14864,II14833
	,II14802,II14771,II14740,II14709,II14678,II14647,II14616,II14585
	,II14554,II14523,II14492,II14461,II14430,II14399,II14368,II14337
	,II14306,II14275,II14244,II14213,II14182,II14151,II14120,II14089
	,II14058,II14027,II10983,II10952,II10921,II10890,II10859,II10828
	,II10797,II10766,II10735,II10704,II10673,II10642,II10611,II10580
	,II10549,II10518,II10487,II10456,II10425,II10394,II10363,II10332
	,II10301,II10270,II10239,II10208,II10177,II10146,II10115,II10084
	,II10053,II10022,II6978,II6947,II6916,II6885,II6854,II6823
	,II6792,II6761,II6730,II6699,II6668,II6637,II6606,II6575
	,II6544,II6513,II6482,II6451,II6420,II6389,II6358,II6327
	,II6296,II6265,II6234,II6203,II6172,II6141,II6110,II6079
	,II6048,II6017,II2973,II2942,II2911,II2880,II2849,II2818
	,II2787,II2756,II2725,II2694,II2663,II2632,II2601,II2570
	,II2539,II2508,II2477,II2446,II2415,II2384,II2353,II2322
	,II2291,II2260,II2229,II2198,II2167,II2136,II2105,II2074
	,II2043,II2012,WX11275,WX11274,WX11273,WX11272,WX11271,WX11270
	,WX11269,WX11268,WX11267,WX11266,WX11265,WX11264,WX11263,WX11262
	,WX11261,WX11260,WX11259,WX11258,WX11257,WX11256,WX11255,WX11254
	,WX11253,WX11252,WX11251,WX11250,WX11249,WX11248,WX11247,WX11246
	,WX11245,WX11244,WX9982,WX9981,WX9980,WX9979,WX9978,WX9977
	,WX9976,WX9975,WX9974,WX9973,WX9972,WX9971,WX9970,WX9969
	,WX9968,WX9967,WX9966,WX9965,WX9964,WX9963,WX9962,WX9961
	,WX9960,WX9959,WX9958,WX9957,WX9956,WX9955,WX9954,WX9953
	,WX9952,WX9951,WX8689,WX8688,WX8687,WX8686,WX8685,WX8684
	,WX8683,WX8682,WX8681,WX8680,WX8679,WX8678,WX8677,WX8676
	,WX8675,WX8674,WX8673,WX8672,WX8671,WX8670,WX8669,WX8668
	,WX8667,WX8666,WX8665,WX8664,WX8663,WX8662,WX8661,WX8660
	,WX8659,WX8658,WX7396,WX7395,WX7394,WX7393,WX7392,WX7391
	,WX7390,WX7389,WX7388,WX7387,WX7386,WX7385,WX7384,WX7383
	,WX7382,WX7381,WX7380,WX7379,WX7378,WX7377,WX7376,WX7375
	,WX7374,WX7373,WX7372,WX7371,WX7370,WX7369,WX7368,WX7367
	,WX7366,WX7365,WX6103,WX6102,WX6101,WX6100,WX6099,WX6098
	,WX6097,WX6096,WX6095,WX6094,WX6093,WX6092,WX6091,WX6090
	,WX6089,WX6088,WX6087,WX6086,WX6085,WX6084,WX6083,WX6082
	,WX6081,WX6080,WX6079,WX6078,WX6077,WX6076,WX6075,WX6074
	,WX6073,WX6072,WX4810,WX4809,WX4808,WX4807,WX4806,WX4805
	,WX4804,WX4803,WX4802,WX4801,WX4800,WX4799,WX4798,WX4797
	,WX4796,WX4795,WX4794,WX4793,WX4792,WX4791,WX4790,WX4789
	,WX4788,WX4787,WX4786,WX4785,WX4784,WX4783,WX4782,WX4781
	,WX4780,WX4779,WX3517,WX3516,WX3515,WX3514,WX3513,WX3512
	,WX3511,WX3510,WX3509,WX3508,WX3507,WX3506,WX3505,WX3504
	,WX3503,WX3502,WX3501,WX3500,WX3499,WX3498,WX3497,WX3496
	,WX3495,WX3494,WX3493,WX3492,WX3491,WX3490,WX3489,WX3488
	,WX3487,WX3486,WX2224,WX2223,WX2222,WX2221,WX2220,WX2219
	,WX2218,WX2217,WX2216,WX2215,WX2214,WX2213,WX2212,WX2211
	,WX2210,WX2209,WX2208,WX2207,WX2206,WX2205,WX2204,WX2203
	,WX2202,WX2201,WX2200,WX2199,WX2198,WX2197,WX2196,WX2195
	,WX2194,WX2193,WX931,WX930,WX929,WX928,WX927,WX926
	,WX925,WX924,WX923,WX922,WX921,WX920,WX919,WX918
	,WX917,WX916,WX915,WX914,WX913,WX912,WX911,WX910
	,WX909,WX908,WX907,WX906,WX905,WX904,WX903,WX902
	,WX901,WX900,WX964,WX966,WX968,WX970,WX972,WX974
	,WX976,WX978,WX980,WX982,WX984,WX986,WX988,WX990
	,WX992,WX994,WX932,WX934,WX936,WX938,WX940,WX942
	,WX944,WX946,WX948,WX950,WX952,WX954,WX956,WX958
	,WX960,WX962,WX2257,WX2259,WX2261,WX2263,WX2265,WX2267
	,WX2269,WX2271,WX2273,WX2275,WX2277,WX2279,WX2281,WX2283
	,WX2285,WX2287,WX2225,WX2227,WX2229,WX2231,WX2233,WX2235
	,WX2237,WX2239,WX2241,WX2243,WX2245,WX2247,WX2249,WX2251
	,WX2253,WX2255,WX3550,WX3552,WX3554,WX3556,WX3558,WX3560
	,WX3562,WX3564,WX3566,WX3568,WX3570,WX3572,WX3574,WX3576
	,WX3578,WX3580,WX3518,WX3520,WX3522,WX3524,WX3526,WX3528
	,WX3530,WX3532,WX3534,WX3536,WX3538,WX3540,WX3542,WX3544
	,WX3546,WX3548,WX4843,WX4845,WX4847,WX4849,WX4851,WX4853
	,WX4855,WX4857,WX4859,WX4861,WX4863,WX4865,WX4867,WX4869
	,WX4871,WX4873,WX4811,WX4813,WX4815,WX4817,WX4819,WX4821
	,WX4823,WX4825,WX4827,WX4829,WX4831,WX4833,WX4835,WX4837
	,WX4839,WX4841,WX6136,WX6138,WX6140,WX6142,WX6144,WX6146
	,WX6148,WX6150,WX6152,WX6154,WX6156,WX6158,WX6160,WX6162
	,WX6164,WX6166,WX6104,WX6106,WX6108,WX6110,WX6112,WX6114
	,WX6116,WX6118,WX6120,WX6122,WX6124,WX6126,WX6128,WX6130
	,WX6132,WX6134,WX7429,WX7431,WX7433,WX7435,WX7437,WX7439
	,WX7441,WX7443,WX7445,WX7447,WX7449,WX7451,WX7453,WX7455
	,WX7457,WX7459,WX7397,WX7399,WX7401,WX7403,WX7405,WX7407
	,WX7409,WX7411,WX7413,WX7415,WX7417,WX7419,WX7421,WX7423
	,WX7425,WX7427,WX8722,WX8724,WX8726,WX8728,WX8730,WX8732
	,WX8734,WX8736,WX8738,WX8740,WX8742,WX8744,WX8746,WX8748
	,WX8750,WX8752,WX8690,WX8692,WX8694,WX8696,WX8698,WX8700
	,WX8702,WX8704,WX8706,WX8708,WX8710,WX8712,WX8714,WX8716
	,WX8718,WX8720,WX10015,WX10017,WX10019,WX10021,WX10023,WX10025
	,WX10027,WX10029,WX10031,WX10033,WX10035,WX10037,WX10039,WX10041
	,WX10043,WX10045,WX9983,WX9985,WX9987,WX9989,WX9991,WX9993
	,WX9995,WX9997,WX9999,WX10001,WX10003,WX10005,WX10007,WX10009
	,WX10011,WX10013,WX11308,WX11310,WX11312,WX11314,WX11316,WX11318
	,WX11320,WX11322,WX11324,WX11326,WX11328,WX11330,WX11332,WX11334
	,WX11336,WX11338,WX11276,WX11278,WX11280,WX11282,WX11284,WX11286
	,WX11288,WX11290,WX11292,WX11294,WX11296,WX11298,WX11300,WX11302
	,WX11304,WX11306,WX11307,WX11305,WX11303,WX11301,WX11299,WX11297
	,WX11295,WX11293,WX11291,WX11289,WX11287,WX11285,WX11283,WX11281
	,WX11279,WX11277,WX11339,WX11337,WX11335,WX11333,WX11331,WX11329
	,WX11327,WX11325,WX11323,WX11321,WX11319,WX11317,WX11315,WX11313
	,WX11311,WX11309,WX10014,WX10012,WX10010,WX10008,WX10006,WX10004
	,WX10002,WX10000,WX9998,WX9996,WX9994,WX9992,WX9990,WX9988
	,WX9986,WX9984,WX10046,WX10044,WX10042,WX10040,WX10038,WX10036
	,WX10034,WX10032,WX10030,WX10028,WX10026,WX10024,WX10022,WX10020
	,WX10018,WX10016,WX8721,WX8719,WX8717,WX8715,WX8713,WX8711
	,WX8709,WX8707,WX8705,WX8703,WX8701,WX8699,WX8697,WX8695
	,WX8693,WX8691,WX8753,WX8751,WX8749,WX8747,WX8745,WX8743
	,WX8741,WX8739,WX8737,WX8735,WX8733,WX8731,WX8729,WX8727
	,WX8725,WX8723,WX7428,WX7426,WX7424,WX7422,WX7420,WX7418
	,WX7416,WX7414,WX7412,WX7410,WX7408,WX7406,WX7404,WX7402
	,WX7400,WX7398,WX7460,WX7458,WX7456,WX7454,WX7452,WX7450
	,WX7448,WX7446,WX7444,WX7442,WX7440,WX7438,WX7436,WX7434
	,WX7432,WX7430,WX6135,WX6133,WX6131,WX6129,WX6127,WX6125
	,WX6123,WX6121,WX6119,WX6117,WX6115,WX6113,WX6111,WX6109
	,WX6107,WX6105,WX6167,WX6165,WX6163,WX6161,WX6159,WX6157
	,WX6155,WX6153,WX6151,WX6149,WX6147,WX6145,WX6143,WX6141
	,WX6139,WX6137,WX4842,WX4840,WX4838,WX4836,WX4834,WX4832
	,WX4830,WX4828,WX4826,WX4824,WX4822,WX4820,WX4818,WX4816
	,WX4814,WX4812,WX4874,WX4872,WX4870,WX4868,WX4866,WX4864
	,WX4862,WX4860,WX4858,WX4856,WX4854,WX4852,WX4850,WX4848
	,WX4846,WX4844,WX3549,WX3547,WX3545,WX3543,WX3541,WX3539
	,WX3537,WX3535,WX3533,WX3531,WX3529,WX3527,WX3525,WX3523
	,WX3521,WX3519,WX3581,WX3579,WX3577,WX3575,WX3573,WX3571
	,WX3569,WX3567,WX3565,WX3563,WX3561,WX3559,WX3557,WX3555
	,WX3553,WX3551,WX2256,WX2254,WX2252,WX2250,WX2248,WX2246
	,WX2244,WX2242,WX2240,WX2238,WX2236,WX2234,WX2232,WX2230
	,WX2228,WX2226,WX2288,WX2286,WX2284,WX2282,WX2280,WX2278
	,WX2276,WX2274,WX2272,WX2270,WX2268,WX2266,WX2264,WX2262
	,WX2260,WX2258,WX963,WX961,WX959,WX957,WX955,WX953
	,WX951,WX949,WX947,WX945,WX943,WX941,WX939,WX937
	,WX935,WX933,WX995,WX993,WX991,WX989,WX987,WX985
	,WX983,WX981,WX979,WX977,WX975,WX973,WX971,WX969
	,WX967,WX965,WX548,WX549,WX550,WX551,WX552,WX553
	,WX554,WX555,WX556,WX557,WX558,WX559,WX560,WX561
	,WX562,WX563,WX564,WX565,WX566,WX567,WX568,WX569
	,WX570,WX571,WX572,WX573,WX574,WX575,WX576,WX577
	,WX578,WX579,WX1841,WX1842,WX1843,WX1844,WX1845,WX1846
	,WX1847,WX1848,WX1849,WX1850,WX1851,WX1852,WX1853,WX1854
	,WX1855,WX1856,WX1857,WX1858,WX1859,WX1860,WX1861,WX1862
	,WX1863,WX1864,WX1865,WX1866,WX1867,WX1868,WX1869,WX1870
	,WX1871,WX1872,WX3134,WX3135,WX3136,WX3137,WX3138,WX3139
	,WX3140,WX3141,WX3142,WX3143,WX3144,WX3145,WX3146,WX3147
	,WX3148,WX3149,WX3150,WX3151,WX3152,WX3153,WX3154,WX3155
	,WX3156,WX3157,WX3158,WX3159,WX3160,WX3161,WX3162,WX3163
	,WX3164,WX3165,WX4427,WX4428,WX4429,WX4430,WX4431,WX4432
	,WX4433,WX4434,WX4435,WX4436,WX4437,WX4438,WX4439,WX4440
	,WX4441,WX4442,WX4443,WX4444,WX4445,WX4446,WX4447,WX4448
	,WX4449,WX4450,WX4451,WX4452,WX4453,WX4454,WX4455,WX4456
	,WX4457,WX4458,WX5720,WX5721,WX5722,WX5723,WX5724,WX5725
	,WX5726,WX5727,WX5728,WX5729,WX5730,WX5731,WX5732,WX5733
	,WX5734,WX5735,WX5736,WX5737,WX5738,WX5739,WX5740,WX5741
	,WX5742,WX5743,WX5744,WX5745,WX5746,WX5747,WX5748,WX5749
	,WX5750,WX5751,WX7013,WX7014,WX7015,WX7016,WX7017,WX7018
	,WX7019,WX7020,WX7021,WX7022,WX7023,WX7024,WX7025,WX7026
	,WX7027,WX7028,WX7029,WX7030,WX7031,WX7032,WX7033,WX7034
	,WX7035,WX7036,WX7037,WX7038,WX7039,WX7040,WX7041,WX7042
	,WX7043,WX7044,WX8306,WX8307,WX8308,WX8309,WX8310,WX8311
	,WX8312,WX8313,WX8314,WX8315,WX8316,WX8317,WX8318,WX8319
	,WX8320,WX8321,WX8322,WX8323,WX8324,WX8325,WX8326,WX8327
	,WX8328,WX8329,WX8330,WX8331,WX8332,WX8333,WX8334,WX8335
	,WX8336,WX8337,WX9599,WX9600,WX9601,WX9602,WX9603,WX9604
	,WX9605,WX9606,WX9607,WX9608,WX9609,WX9610,WX9611,WX9612
	,WX9613,WX9614,WX9615,WX9616,WX9617,WX9618,WX9619,WX9620
	,WX9621,WX9622,WX9623,WX9624,WX9625,WX9626,WX9627,WX9628
	,WX9629,WX9630,WX10892,WX10893,WX10894,WX10895,WX10896,WX10897
	,WX10898,WX10899,WX10900,WX10901,WX10902,WX10903,WX10904,WX10905
	,WX10906,WX10907,WX10908,WX10909,WX10910,WX10911,WX10912,WX10913
	,WX10914,WX10915,WX10916,WX10917,WX10918,WX10919,WX10920,WX10921
	,WX10922,WX10923,WX10955,WX10954,WX10953,WX10952,WX10951,WX10950
	,WX10949,WX10948,WX10947,WX10946,WX10945,WX10944,WX10943,WX10942
	,WX10941,WX10940,WX10939,WX10938,WX10937,WX10936,WX10935,WX10934
	,WX10933,WX10932,WX10931,WX10930,WX10929,WX10928,WX10927,WX10926
	,WX10925,WX10924,WX9662,WX9661,WX9660,WX9659,WX9658,WX9657
	,WX9656,WX9655,WX9654,WX9653,WX9652,WX9651,WX9650,WX9649
	,WX9648,WX9647,WX9646,WX9645,WX9644,WX9643,WX9642,WX9641
	,WX9640,WX9639,WX9638,WX9637,WX9636,WX9635,WX9634,WX9633
	,WX9632,WX9631,WX8369,WX8368,WX8367,WX8366,WX8365,WX8364
	,WX8363,WX8362,WX8361,WX8360,WX8359,WX8358,WX8357,WX8356
	,WX8355,WX8354,WX8353,WX8352,WX8351,WX8350,WX8349,WX8348
	,WX8347,WX8346,WX8345,WX8344,WX8343,WX8342,WX8341,WX8340
	,WX8339,WX8338,WX7076,WX7075,WX7074,WX7073,WX7072,WX7071
	,WX7070,WX7069,WX7068,WX7067,WX7066,WX7065,WX7064,WX7063
	,WX7062,WX7061,WX7060,WX7059,WX7058,WX7057,WX7056,WX7055
	,WX7054,WX7053,WX7052,WX7051,WX7050,WX7049,WX7048,WX7047
	,WX7046,WX7045,WX5783,WX5782,WX5781,WX5780,WX5779,WX5778
	,WX5777,WX5776,WX5775,WX5774,WX5773,WX5772,WX5771,WX5770
	,WX5769,WX5768,WX5767,WX5766,WX5765,WX5764,WX5763,WX5762
	,WX5761,WX5760,WX5759,WX5758,WX5757,WX5756,WX5755,WX5754
	,WX5753,WX5752,WX4490,WX4489,WX4488,WX4487,WX4486,WX4485
	,WX4484,WX4483,WX4482,WX4481,WX4480,WX4479,WX4478,WX4477
	,WX4476,WX4475,WX4474,WX4473,WX4472,WX4471,WX4470,WX4469
	,WX4468,WX4467,WX4466,WX4465,WX4464,WX4463,WX4462,WX4461
	,WX4460,WX4459,WX3197,WX3196,WX3195,WX3194,WX3193,WX3192
	,WX3191,WX3190,WX3189,WX3188,WX3187,WX3186,WX3185,WX3184
	,WX3183,WX3182,WX3181,WX3180,WX3179,WX3178,WX3177,WX3176
	,WX3175,WX3174,WX3173,WX3172,WX3171,WX3170,WX3169,WX3168
	,WX3167,WX3166,WX1904,WX1903,WX1902,WX1901,WX1900,WX1899
	,WX1898,WX1897,WX1896,WX1895,WX1894,WX1893,WX1892,WX1891
	,WX1890,WX1889,WX1888,WX1887,WX1886,WX1885,WX1884,WX1883
	,WX1882,WX1881,WX1880,WX1879,WX1878,WX1877,WX1876,WX1875
	,WX1874,WX1873,WX611,WX610,WX609,WX608,WX607,WX606
	,WX605,WX604,WX603,WX602,WX601,WX600,WX599,WX598
	,WX597,WX596,WX595,WX594,WX593,WX592,WX591,WX590
	,WX589,WX588,WX587,WX586,WX585,WX584,WX583,WX582
	,WX581,WX580,WX11569,WX11562,WX11555,WX11548,WX11541,WX11534
	,WX11527,WX11520,WX11513,WX11506,WX11499,WX11492,WX11485,WX11478
	,WX11471,WX11464,WX11457,WX11450,WX11443,WX11436,WX11429,WX11422
	,WX11415,WX11408,WX11401,WX11394,WX11387,WX11380,WX11373,WX11366
	,WX11359,WX11352,WX10276,WX10269,WX10262,WX10255,WX10248,WX10241
	,WX10234,WX10227,WX10220,WX10213,WX10206,WX10199,WX10192,WX10185
	,WX10178,WX10171,WX10164,WX10157,WX10150,WX10143,WX10136,WX10129
	,WX10122,WX10115,WX10108,WX10101,WX10094,WX10087,WX10080,WX10073
	,WX10066,WX10059,WX8983,WX8976,WX8969,WX8962,WX8955,WX8948
	,WX8941,WX8934,WX8927,WX8920,WX8913,WX8906,WX8899,WX8892
	,WX8885,WX8878,WX8871,WX8864,WX8857,WX8850,WX8843,WX8836
	,WX8829,WX8822,WX8815,WX8808,WX8801,WX8794,WX8787,WX8780
	,WX8773,WX8766,WX7690,WX7683,WX7676,WX7669,WX7662,WX7655
	,WX7648,WX7641,WX7634,WX7627,WX7620,WX7613,WX7606,WX7599
	,WX7592,WX7585,WX7578,WX7571,WX7564,WX7557,WX7550,WX7543
	,WX7536,WX7529,WX7522,WX7515,WX7508,WX7501,WX7494,WX7487
	,WX7480,WX7473,WX6397,WX6390,WX6383,WX6376,WX6369,WX6362
	,WX6355,WX6348,WX6341,WX6334,WX6327,WX6320,WX6313,WX6306
	,WX6299,WX6292,WX6285,WX6278,WX6271,WX6264,WX6257,WX6250
	,WX6243,WX6236,WX6229,WX6222,WX6215,WX6208,WX6201,WX6194
	,WX6187,WX6180,WX5104,WX5097,WX5090,WX5083,WX5076,WX5069
	,WX5062,WX5055,WX5048,WX5041,WX5034,WX5027,WX5020,WX5013
	,WX5006,WX4999,WX4992,WX4985,WX4978,WX4971,WX4964,WX4957
	,WX4950,WX4943,WX4936,WX4929,WX4922,WX4915,WX4908,WX4901
	,WX4894,WX4887,WX3811,WX3804,WX3797,WX3790,WX3783,WX3776
	,WX3769,WX3762,WX3755,WX3748,WX3741,WX3734,WX3727,WX3720
	,WX3713,WX3706,WX3699,WX3692,WX3685,WX3678,WX3671,WX3664
	,WX3657,WX3650,WX3643,WX3636,WX3629,WX3622,WX3615,WX3608
	,WX3601,WX3594,WX2518,WX2511,WX2504,WX2497,WX2490,WX2483
	,WX2476,WX2469,WX2462,WX2455,WX2448,WX2441,WX2434,WX2427
	,WX2420,WX2413,WX2406,WX2399,WX2392,WX2385,WX2378,WX2371
	,WX2364,WX2357,WX2350,WX2343,WX2336,WX2329,WX2322,WX2315
	,WX2308,WX2301,WX1225,WX1218,WX1211,WX1204,WX1197,WX1190
	,WX1183,WX1176,WX1169,WX1162,WX1155,WX1148,WX1141,WX1134
	,WX1127,WX1120,WX1113,WX1106,WX1099,WX1092,WX1085,WX1078
	,WX1071,WX1064,WX1057,WX1050,WX1043,WX1036,WX1029,WX1022
	,WX1015,WX1008,II3052,II3065,II3078,II3091,II3104,II3117
	,II3130,II3143,II3156,II3169,II3182,II3195,II3208,II3221
	,II3234,II3247,II3260,II3273,II3286,II3299,II3312,II3325
	,II3338,II3351,II3364,II3377,II3390,II3403,II3416,II3429
	,II3442,II3455,II7057,II7070,II7083,II7096,II7109,II7122
	,II7135,II7148,II7161,II7174,II7187,II7200,II7213,II7226
	,II7239,II7252,II7265,II7278,II7291,II7304,II7317,II7330
	,II7343,II7356,II7369,II7382,II7395,II7408,II7421,II7434
	,II7447,II7460,II11062,II11075,II11088,II11101,II11114,II11127
	,II11140,II11153,II11166,II11179,II11192,II11205,II11218,II11231
	,II11244,II11257,II11270,II11283,II11296,II11309,II11322,II11335
	,II11348,II11361,II11374,II11387,II11400,II11413,II11426,II11439
	,II11452,II11465,II15067,II15080,II15093,II15106,II15119,II15132
	,II15145,II15158,II15171,II15184,II15197,II15210,II15223,II15236
	,II15249,II15262,II15275,II15288,II15301,II15314,II15327,II15340
	,II15353,II15366,II15379,II15392,II15405,II15418,II15431,II15444
	,II15457,II15470,II19072,II19085,II19098,II19111,II19124,II19137
	,II19150,II19163,II19176,II19189,II19202,II19215,II19228,II19241
	,II19254,II19267,II19280,II19293,II19306,II19319,II19332,II19345
	,II19358,II19371,II19384,II19397,II19410,II19423,II19436,II19449
	,II19462,II19475,II23077,II23090,II23103,II23116,II23129,II23142
	,II23155,II23168,II23181,II23194,II23207,II23220,II23233,II23246
	,II23259,II23272,II23285,II23298,II23311,II23324,II23337,II23350
	,II23363,II23376,II23389,II23402,II23415,II23428,II23441,II23454
	,II23467,II23480,II27082,II27095,II27108,II27121,II27134,II27147
	,II27160,II27173,II27186,II27199,II27212,II27225,II27238,II27251
	,II27264,II27277,II27290,II27303,II27316,II27329,II27342,II27355
	,II27368,II27381,II27394,II27407,II27420,II27433,II27446,II27459
	,II27472,II27485,II31087,II31100,II31113,II31126,II31139,II31152
	,II31165,II31178,II31191,II31204,II31217,II31230,II31243,II31256
	,II31269,II31282,II31295,II31308,II31321,II31334,II31347,II31360
	,II31373,II31386,II31399,II31412,II31425,II31438,II31451,II31464
	,II31477,II31490,II35092,II35105,II35118,II35131,II35144,II35157
	,II35170,II35183,II35196,II35209,II35222,II35235,II35248,II35261
	,II35274,II35287,II35300,II35313,II35326,II35339,II35352,II35365
	,II35378,II35391,II35404,II35417,II35430,II35443,II35456,II35469
	,II35482,II35495,II35496,II35483,II35470,II35457,II35444,II35431
	,II35418,II35405,II35392,II35379,II35366,II35353,II35340,II35327
	,II35314,II35301,II35288,II35275,II35262,II35249,II35236,II35223
	,II35210,II35197,II35184,II35171,II35158,II35145,II35132,II35119
	,II35106,II35093,II31491,II31478,II31465,II31452,II31439,II31426
	,II31413,II31400,II31387,II31374,II31361,II31348,II31335,II31322
	,II31309,II31296,II31283,II31270,II31257,II31244,II31231,II31218
	,II31205,II31192,II31179,II31166,II31153,II31140,II31127,II31114
	,II31101,II31088,II27486,II27473,II27460,II27447,II27434,II27421
	,II27408,II27395,II27382,II27369,II27356,II27343,II27330,II27317
	,II27304,II27291,II27278,II27265,II27252,II27239,II27226,II27213
	,II27200,II27187,II27174,II27161,II27148,II27135,II27122,II27109
	,II27096,II27083,II23481,II23468,II23455,II23442,II23429,II23416
	,II23403,II23390,II23377,II23364,II23351,II23338,II23325,II23312
	,II23299,II23286,II23273,II23260,II23247,II23234,II23221,II23208
	,II23195,II23182,II23169,II23156,II23143,II23130,II23117,II23104
	,II23091,II23078,II19476,II19463,II19450,II19437,II19424,II19411
	,II19398,II19385,II19372,II19359,II19346,II19333,II19320,II19307
	,II19294,II19281,II19268,II19255,II19242,II19229,II19216,II19203
	,II19190,II19177,II19164,II19151,II19138,II19125,II19112,II19099
	,II19086,II19073,II15471,II15458,II15445,II15432,II15419,II15406
	,II15393,II15380,II15367,II15354,II15341,II15328,II15315,II15302
	,II15289,II15276,II15263,II15250,II15237,II15224,II15211,II15198
	,II15185,II15172,II15159,II15146,II15133,II15120,II15107,II15094
	,II15081,II15068,II11466,II11453,II11440,II11427,II11414,II11401
	,II11388,II11375,II11362,II11349,II11336,II11323,II11310,II11297
	,II11284,II11271,II11258,II11245,II11232,II11219,II11206,II11193
	,II11180,II11167,II11154,II11141,II11128,II11115,II11102,II11089
	,II11076,II11063,II7461,II7448,II7435,II7422,II7409,II7396
	,II7383,II7370,II7357,II7344,II7331,II7318,II7305,II7292
	,II7279,II7266,II7253,II7240,II7227,II7214,II7201,II7188
	,II7175,II7162,II7149,II7136,II7123,II7110,II7097,II7084
	,II7071,II7058,II3456,II3443,II3430,II3417,II3404,II3391
	,II3378,II3365,II3352,II3339,II3326,II3313,II3300,II3287
	,II3274,II3261,II3248,II3235,II3222,II3209,II3196,II3183
	,II3170,II3157,II3144,II3131,II3118,II3105,II3092,II3079
	,II3066,II3053,II3054,II3067,II3080,II3093,II3106,II3119
	,II3132,II3145,II3158,II3171,II3184,II3197,II3210,II3223
	,II3236,II3249,II3262,II3275,II3288,II3301,II3314,II3327
	,II3340,II3353,II3366,II3379,II3392,II3405,II3418,II3431
	,II3444,II3457,II7059,II7072,II7085,II7098,II7111,II7124
	,II7137,II7150,II7163,II7176,II7189,II7202,II7215,II7228
	,II7241,II7254,II7267,II7280,II7293,II7306,II7319,II7332
	,II7345,II7358,II7371,II7384,II7397,II7410,II7423,II7436
	,II7449,II7462,II11064,II11077,II11090,II11103,II11116,II11129
	,II11142,II11155,II11168,II11181,II11194,II11207,II11220,II11233
	,II11246,II11259,II11272,II11285,II11298,II11311,II11324,II11337
	,II11350,II11363,II11376,II11389,II11402,II11415,II11428,II11441
	,II11454,II11467,II15069,II15082,II15095,II15108,II15121,II15134
	,II15147,II15160,II15173,II15186,II15199,II15212,II15225,II15238
	,II15251,II15264,II15277,II15290,II15303,II15316,II15329,II15342
	,II15355,II15368,II15381,II15394,II15407,II15420,II15433,II15446
	,II15459,II15472,II19074,II19087,II19100,II19113,II19126,II19139
	,II19152,II19165,II19178,II19191,II19204,II19217,II19230,II19243
	,II19256,II19269,II19282,II19295,II19308,II19321,II19334,II19347
	,II19360,II19373,II19386,II19399,II19412,II19425,II19438,II19451
	,II19464,II19477,II23079,II23092,II23105,II23118,II23131,II23144
	,II23157,II23170,II23183,II23196,II23209,II23222,II23235,II23248
	,II23261,II23274,II23287,II23300,II23313,II23326,II23339,II23352
	,II23365,II23378,II23391,II23404,II23417,II23430,II23443,II23456
	,II23469,II23482,II27084,II27097,II27110,II27123,II27136,II27149
	,II27162,II27175,II27188,II27201,II27214,II27227,II27240,II27253
	,II27266,II27279,II27292,II27305,II27318,II27331,II27344,II27357
	,II27370,II27383,II27396,II27409,II27422,II27435,II27448,II27461
	,II27474,II27487,II31089,II31102,II31115,II31128,II31141,II31154
	,II31167,II31180,II31193,II31206,II31219,II31232,II31245,II31258
	,II31271,II31284,II31297,II31310,II31323,II31336,II31349,II31362
	,II31375,II31388,II31401,II31414,II31427,II31440,II31453,II31466
	,II31479,II31492,II35094,II35107,II35120,II35133,II35146,II35159
	,II35172,II35185,II35198,II35211,II35224,II35237,II35250,II35263
	,II35276,II35289,II35302,II35315,II35328,II35341,II35354,II35367
	,II35380,II35393,II35406,II35419,II35432,II35445,II35458,II35471
	,II35484,II35497,WX1006,WX1013,WX1020,WX1027,WX1034,WX1041
	,WX1048,WX1055,WX1062,WX1069,WX1076,WX1083,WX1090,WX1097
	,WX1104,WX1111,WX1118,WX1125,WX1132,WX1139,WX1146,WX1153
	,WX1160,WX1167,WX1174,WX1181,WX1188,WX1195,WX1202,WX1209
	,WX1216,WX1223,WX2299,WX2306,WX2313,WX2320,WX2327,WX2334
	,WX2341,WX2348,WX2355,WX2362,WX2369,WX2376,WX2383,WX2390
	,WX2397,WX2404,WX2411,WX2418,WX2425,WX2432,WX2439,WX2446
	,WX2453,WX2460,WX2467,WX2474,WX2481,WX2488,WX2495,WX2502
	,WX2509,WX2516,WX3592,WX3599,WX3606,WX3613,WX3620,WX3627
	,WX3634,WX3641,WX3648,WX3655,WX3662,WX3669,WX3676,WX3683
	,WX3690,WX3697,WX3704,WX3711,WX3718,WX3725,WX3732,WX3739
	,WX3746,WX3753,WX3760,WX3767,WX3774,WX3781,WX3788,WX3795
	,WX3802,WX3809,WX4885,WX4892,WX4899,WX4906,WX4913,WX4920
	,WX4927,WX4934,WX4941,WX4948,WX4955,WX4962,WX4969,WX4976
	,WX4983,WX4990,WX4997,WX5004,WX5011,WX5018,WX5025,WX5032
	,WX5039,WX5046,WX5053,WX5060,WX5067,WX5074,WX5081,WX5088
	,WX5095,WX5102,WX6178,WX6185,WX6192,WX6199,WX6206,WX6213
	,WX6220,WX6227,WX6234,WX6241,WX6248,WX6255,WX6262,WX6269
	,WX6276,WX6283,WX6290,WX6297,WX6304,WX6311,WX6318,WX6325
	,WX6332,WX6339,WX6346,WX6353,WX6360,WX6367,WX6374,WX6381
	,WX6388,WX6395,WX7471,WX7478,WX7485,WX7492,WX7499,WX7506
	,WX7513,WX7520,WX7527,WX7534,WX7541,WX7548,WX7555,WX7562
	,WX7569,WX7576,WX7583,WX7590,WX7597,WX7604,WX7611,WX7618
	,WX7625,WX7632,WX7639,WX7646,WX7653,WX7660,WX7667,WX7674
	,WX7681,WX7688,WX8764,WX8771,WX8778,WX8785,WX8792,WX8799
	,WX8806,WX8813,WX8820,WX8827,WX8834,WX8841,WX8848,WX8855
	,WX8862,WX8869,WX8876,WX8883,WX8890,WX8897,WX8904,WX8911
	,WX8918,WX8925,WX8932,WX8939,WX8946,WX8953,WX8960,WX8967
	,WX8974,WX8981,WX10057,WX10064,WX10071,WX10078,WX10085,WX10092
	,WX10099,WX10106,WX10113,WX10120,WX10127,WX10134,WX10141,WX10148
	,WX10155,WX10162,WX10169,WX10176,WX10183,WX10190,WX10197,WX10204
	,WX10211,WX10218,WX10225,WX10232,WX10239,WX10246,WX10253,WX10260
	,WX10267,WX10274,WX11350,WX11357,WX11364,WX11371,WX11378,WX11385
	,WX11392,WX11399,WX11406,WX11413,WX11420,WX11427,WX11434,WX11441
	,WX11448,WX11455,WX11462,WX11469,WX11476,WX11483,WX11490,WX11497
	,WX11504,WX11511,WX11518,WX11525,WX11532,WX11539,WX11546,WX11553
	,WX11560,WX11567,WX11568,WX11561,WX11554,WX11547,WX11540,WX11533
	,WX11526,WX11519,WX11512,WX11505,WX11498,WX11491,WX11484,WX11477
	,WX11470,WX11463,WX11456,WX11449,WX11442,WX11435,WX11428,WX11421
	,WX11414,WX11407,WX11400,WX11393,WX11386,WX11379,WX11372,WX11365
	,WX11358,WX11351,WX10275,WX10268,WX10261,WX10254,WX10247,WX10240
	,WX10233,WX10226,WX10219,WX10212,WX10205,WX10198,WX10191,WX10184
	,WX10177,WX10170,WX10163,WX10156,WX10149,WX10142,WX10135,WX10128
	,WX10121,WX10114,WX10107,WX10100,WX10093,WX10086,WX10079,WX10072
	,WX10065,WX10058,WX8982,WX8975,WX8968,WX8961,WX8954,WX8947
	,WX8940,WX8933,WX8926,WX8919,WX8912,WX8905,WX8898,WX8891
	,WX8884,WX8877,WX8870,WX8863,WX8856,WX8849,WX8842,WX8835
	,WX8828,WX8821,WX8814,WX8807,WX8800,WX8793,WX8786,WX8779
	,WX8772,WX8765,WX7689,WX7682,WX7675,WX7668,WX7661,WX7654
	,WX7647,WX7640,WX7633,WX7626,WX7619,WX7612,WX7605,WX7598
	,WX7591,WX7584,WX7577,WX7570,WX7563,WX7556,WX7549,WX7542
	,WX7535,WX7528,WX7521,WX7514,WX7507,WX7500,WX7493,WX7486
	,WX7479,WX7472,WX6396,WX6389,WX6382,WX6375,WX6368,WX6361
	,WX6354,WX6347,WX6340,WX6333,WX6326,WX6319,WX6312,WX6305
	,WX6298,WX6291,WX6284,WX6277,WX6270,WX6263,WX6256,WX6249
	,WX6242,WX6235,WX6228,WX6221,WX6214,WX6207,WX6200,WX6193
	,WX6186,WX6179,WX5103,WX5096,WX5089,WX5082,WX5075,WX5068
	,WX5061,WX5054,WX5047,WX5040,WX5033,WX5026,WX5019,WX5012
	,WX5005,WX4998,WX4991,WX4984,WX4977,WX4970,WX4963,WX4956
	,WX4949,WX4942,WX4935,WX4928,WX4921,WX4914,WX4907,WX4900
	,WX4893,WX4886,WX3810,WX3803,WX3796,WX3789,WX3782,WX3775
	,WX3768,WX3761,WX3754,WX3747,WX3740,WX3733,WX3726,WX3719
	,WX3712,WX3705,WX3698,WX3691,WX3684,WX3677,WX3670,WX3663
	,WX3656,WX3649,WX3642,WX3635,WX3628,WX3621,WX3614,WX3607
	,WX3600,WX3593,WX2517,WX2510,WX2503,WX2496,WX2489,WX2482
	,WX2475,WX2468,WX2461,WX2454,WX2447,WX2440,WX2433,WX2426
	,WX2419,WX2412,WX2405,WX2398,WX2391,WX2384,WX2377,WX2370
	,WX2363,WX2356,WX2349,WX2342,WX2335,WX2328,WX2321,WX2314
	,WX2307,WX2300,WX1224,WX1217,WX1210,WX1203,WX1196,WX1189
	,WX1182,WX1175,WX1168,WX1161,WX1154,WX1147,WX1140,WX1133
	,WX1126,WX1119,WX1112,WX1105,WX1098,WX1091,WX1084,WX1077
	,WX1070,WX1063,WX1056,WX1049,WX1042,WX1035,WX1028,WX1021
	,WX1014,WX1007,WX1010,WX1017,WX1024,WX1031,WX1038,WX1045
	,WX1052,WX1059,WX1066,WX1073,WX1080,WX1087,WX1094,WX1101
	,WX1108,WX1115,WX1122,WX1129,WX1136,WX1143,WX1150,WX1157
	,WX1164,WX1171,WX1178,WX1185,WX1192,WX1199,WX1206,WX1213
	,WX1220,WX1227,WX2303,WX2310,WX2317,WX2324,WX2331,WX2338
	,WX2345,WX2352,WX2359,WX2366,WX2373,WX2380,WX2387,WX2394
	,WX2401,WX2408,WX2415,WX2422,WX2429,WX2436,WX2443,WX2450
	,WX2457,WX2464,WX2471,WX2478,WX2485,WX2492,WX2499,WX2506
	,WX2513,WX2520,WX3596,WX3603,WX3610,WX3617,WX3624,WX3631
	,WX3638,WX3645,WX3652,WX3659,WX3666,WX3673,WX3680,WX3687
	,WX3694,WX3701,WX3708,WX3715,WX3722,WX3729,WX3736,WX3743
	,WX3750,WX3757,WX3764,WX3771,WX3778,WX3785,WX3792,WX3799
	,WX3806,WX3813,WX4889,WX4896,WX4903,WX4910,WX4917,WX4924
	,WX4931,WX4938,WX4945,WX4952,WX4959,WX4966,WX4973,WX4980
	,WX4987,WX4994,WX5001,WX5008,WX5015,WX5022,WX5029,WX5036
	,WX5043,WX5050,WX5057,WX5064,WX5071,WX5078,WX5085,WX5092
	,WX5099,WX5106,WX6182,WX6189,WX6196,WX6203,WX6210,WX6217
	,WX6224,WX6231,WX6238,WX6245,WX6252,WX6259,WX6266,WX6273
	,WX6280,WX6287,WX6294,WX6301,WX6308,WX6315,WX6322,WX6329
	,WX6336,WX6343,WX6350,WX6357,WX6364,WX6371,WX6378,WX6385
	,WX6392,WX6399,WX7475,WX7482,WX7489,WX7496,WX7503,WX7510
	,WX7517,WX7524,WX7531,WX7538,WX7545,WX7552,WX7559,WX7566
	,WX7573,WX7580,WX7587,WX7594,WX7601,WX7608,WX7615,WX7622
	,WX7629,WX7636,WX7643,WX7650,WX7657,WX7664,WX7671,WX7678
	,WX7685,WX7692,WX8768,WX8775,WX8782,WX8789,WX8796,WX8803
	,WX8810,WX8817,WX8824,WX8831,WX8838,WX8845,WX8852,WX8859
	,WX8866,WX8873,WX8880,WX8887,WX8894,WX8901,WX8908,WX8915
	,WX8922,WX8929,WX8936,WX8943,WX8950,WX8957,WX8964,WX8971
	,WX8978,WX8985,WX10061,WX10068,WX10075,WX10082,WX10089,WX10096
	,WX10103,WX10110,WX10117,WX10124,WX10131,WX10138,WX10145,WX10152
	,WX10159,WX10166,WX10173,WX10180,WX10187,WX10194,WX10201,WX10208
	,WX10215,WX10222,WX10229,WX10236,WX10243,WX10250,WX10257,WX10264
	,WX10271,WX10278,WX11354,WX11361,WX11368,WX11375,WX11382,WX11389
	,WX11396,WX11403,WX11410,WX11417,WX11424,WX11431,WX11438,WX11445
	,WX11452,WX11459,WX11466,WX11473,WX11480,WX11487,WX11494,WX11501
	,WX11508,WX11515,WX11522,WX11529,WX11536,WX11543,WX11550,WX11557
	,WX11564,WX11571,WX11572,WX11565,WX11558,WX11551,WX11544,WX11537
	,WX11530,WX11523,WX11516,WX11509,WX11502,WX11495,WX11488,WX11481
	,WX11474,WX11467,WX11460,WX11453,WX11446,WX11439,WX11432,WX11425
	,WX11418,WX11411,WX11404,WX11397,WX11390,WX11383,WX11376,WX11369
	,WX11362,WX11355,WX10279,WX10272,WX10265,WX10258,WX10251,WX10244
	,WX10237,WX10230,WX10223,WX10216,WX10209,WX10202,WX10195,WX10188
	,WX10181,WX10174,WX10167,WX10160,WX10153,WX10146,WX10139,WX10132
	,WX10125,WX10118,WX10111,WX10104,WX10097,WX10090,WX10083,WX10076
	,WX10069,WX10062,WX8986,WX8979,WX8972,WX8965,WX8958,WX8951
	,WX8944,WX8937,WX8930,WX8923,WX8916,WX8909,WX8902,WX8895
	,WX8888,WX8881,WX8874,WX8867,WX8860,WX8853,WX8846,WX8839
	,WX8832,WX8825,WX8818,WX8811,WX8804,WX8797,WX8790,WX8783
	,WX8776,WX8769,WX7693,WX7686,WX7679,WX7672,WX7665,WX7658
	,WX7651,WX7644,WX7637,WX7630,WX7623,WX7616,WX7609,WX7602
	,WX7595,WX7588,WX7581,WX7574,WX7567,WX7560,WX7553,WX7546
	,WX7539,WX7532,WX7525,WX7518,WX7511,WX7504,WX7497,WX7490
	,WX7483,WX7476,WX6400,WX6393,WX6386,WX6379,WX6372,WX6365
	,WX6358,WX6351,WX6344,WX6337,WX6330,WX6323,WX6316,WX6309
	,WX6302,WX6295,WX6288,WX6281,WX6274,WX6267,WX6260,WX6253
	,WX6246,WX6239,WX6232,WX6225,WX6218,WX6211,WX6204,WX6197
	,WX6190,WX6183,WX5107,WX5100,WX5093,WX5086,WX5079,WX5072
	,WX5065,WX5058,WX5051,WX5044,WX5037,WX5030,WX5023,WX5016
	,WX5009,WX5002,WX4995,WX4988,WX4981,WX4974,WX4967,WX4960
	,WX4953,WX4946,WX4939,WX4932,WX4925,WX4918,WX4911,WX4904
	,WX4897,WX4890,WX3814,WX3807,WX3800,WX3793,WX3786,WX3779
	,WX3772,WX3765,WX3758,WX3751,WX3744,WX3737,WX3730,WX3723
	,WX3716,WX3709,WX3702,WX3695,WX3688,WX3681,WX3674,WX3667
	,WX3660,WX3653,WX3646,WX3639,WX3632,WX3625,WX3618,WX3611
	,WX3604,WX3597,WX2521,WX2514,WX2507,WX2500,WX2493,WX2486
	,WX2479,WX2472,WX2465,WX2458,WX2451,WX2444,WX2437,WX2430
	,WX2423,WX2416,WX2409,WX2402,WX2395,WX2388,WX2381,WX2374
	,WX2367,WX2360,WX2353,WX2346,WX2339,WX2332,WX2325,WX2318
	,WX2311,WX2304,WX1228,WX1221,WX1214,WX1207,WX1200,WX1193
	,WX1186,WX1179,WX1172,WX1165,WX1158,WX1151,WX1144,WX1137
	,WX1130,WX1123,WX1116,WX1109,WX1102,WX1095,WX1088,WX1081
	,WX1074,WX1067,WX1060,WX1053,WX1046,WX1039,WX1032,WX1025
	,WX1018,WX1011,WX2305,WX2312,WX2319,WX2326,WX2333,WX2340
	,WX2347,WX2354,WX2361,WX2368,WX2375,WX2382,WX2389,WX2396
	,WX2403,WX2410,WX2417,WX2424,WX2431,WX2438,WX2445,WX2452
	,WX2459,WX2466,WX2473,WX2480,WX2487,WX2494,WX2501,WX2508
	,WX2515,WX2522,WX3598,WX3605,WX3612,WX3619,WX3626,WX3633
	,WX3640,WX3647,WX3654,WX3661,WX3668,WX3675,WX3682,WX3689
	,WX3696,WX3703,WX3710,WX3717,WX3724,WX3731,WX3738,WX3745
	,WX3752,WX3759,WX3766,WX3773,WX3780,WX3787,WX3794,WX3801
	,WX3808,WX3815,WX4891,WX4898,WX4905,WX4912,WX4919,WX4926
	,WX4933,WX4940,WX4947,WX4954,WX4961,WX4968,WX4975,WX4982
	,WX4989,WX4996,WX5003,WX5010,WX5017,WX5024,WX5031,WX5038
	,WX5045,WX5052,WX5059,WX5066,WX5073,WX5080,WX5087,WX5094
	,WX5101,WX5108,WX6184,WX6191,WX6198,WX6205,WX6212,WX6219
	,WX6226,WX6233,WX6240,WX6247,WX6254,WX6261,WX6268,WX6275
	,WX6282,WX6289,WX6296,WX6303,WX6310,WX6317,WX6324,WX6331
	,WX6338,WX6345,WX6352,WX6359,WX6366,WX6373,WX6380,WX6387
	,WX6394,WX6401,WX7477,WX7484,WX7491,WX7498,WX7505,WX7512
	,WX7519,WX7526,WX7533,WX7540,WX7547,WX7554,WX7561,WX7568
	,WX7575,WX7582,WX7589,WX7596,WX7603,WX7610,WX7617,WX7624
	,WX7631,WX7638,WX7645,WX7652,WX7659,WX7666,WX7673,WX7680
	,WX7687,WX7694,WX8770,WX8777,WX8784,WX8791,WX8798,WX8805
	,WX8812,WX8819,WX8826,WX8833,WX8840,WX8847,WX8854,WX8861
	,WX8868,WX8875,WX8882,WX8889,WX8896,WX8903,WX8910,WX8917
	,WX8924,WX8931,WX8938,WX8945,WX8952,WX8959,WX8966,WX8973
	,WX8980,WX8987,WX10063,WX10070,WX10077,WX10084,WX10091,WX10098
	,WX10105,WX10112,WX10119,WX10126,WX10133,WX10140,WX10147,WX10154
	,WX10161,WX10168,WX10175,WX10182,WX10189,WX10196,WX10203,WX10210
	,WX10217,WX10224,WX10231,WX10238,WX10245,WX10252,WX10259,WX10266
	,WX10273,WX10280,WX11356,WX11363,WX11370,WX11377,WX11384,WX11391
	,WX11398,WX11405,WX11412,WX11419,WX11426,WX11433,WX11440,WX11447
	,WX11454,WX11461,WX11468,WX11475,WX11482,WX11489,WX11496,WX11503
	,WX11510,WX11517,WX11524,WX11531,WX11538,WX11545,WX11552,WX11559
	,WX11566,WX11573,WX10822,WX10808,WX10794,WX10780,WX10766,WX10752
	,WX10738,WX10724,WX10710,WX10696,WX10682,WX10668,WX10654,WX10640
	,WX10626,WX10612,WX10598,WX10584,WX10570,WX10556,WX10542,WX10528
	,WX10514,WX10500,WX10486,WX10472,WX10458,WX10444,WX10430,WX10416
	,WX10402,WX10388,WX9529,WX9515,WX9501,WX9487,WX9473,WX9459
	,WX9445,WX9431,WX9417,WX9403,WX9389,WX9375,WX9361,WX9347
	,WX9333,WX9319,WX9305,WX9291,WX9277,WX9263,WX9249,WX9235
	,WX9221,WX9207,WX9193,WX9179,WX9165,WX9151,WX9137,WX9123
	,WX9109,WX9095,WX8236,WX8222,WX8208,WX8194,WX8180,WX8166
	,WX8152,WX8138,WX8124,WX8110,WX8096,WX8082,WX8068,WX8054
	,WX8040,WX8026,WX8012,WX7998,WX7984,WX7970,WX7956,WX7942
	,WX7928,WX7914,WX7900,WX7886,WX7872,WX7858,WX7844,WX7830
	,WX7816,WX7802,WX6943,WX6929,WX6915,WX6901,WX6887,WX6873
	,WX6859,WX6845,WX6831,WX6817,WX6803,WX6789,WX6775,WX6761
	,WX6747,WX6733,WX6719,WX6705,WX6691,WX6677,WX6663,WX6649
	,WX6635,WX6621,WX6607,WX6593,WX6579,WX6565,WX6551,WX6537
	,WX6523,WX6509,WX5650,WX5636,WX5622,WX5608,WX5594,WX5580
	,WX5566,WX5552,WX5538,WX5524,WX5510,WX5496,WX5482,WX5468
	,WX5454,WX5440,WX5426,WX5412,WX5398,WX5384,WX5370,WX5356
	,WX5342,WX5328,WX5314,WX5300,WX5286,WX5272,WX5258,WX5244
	,WX5230,WX5216,WX4357,WX4343,WX4329,WX4315,WX4301,WX4287
	,WX4273,WX4259,WX4245,WX4231,WX4217,WX4203,WX4189,WX4175
	,WX4161,WX4147,WX4133,WX4119,WX4105,WX4091,WX4077,WX4063
	,WX4049,WX4035,WX4021,WX4007,WX3993,WX3979,WX3965,WX3951
	,WX3937,WX3923,WX3064,WX3050,WX3036,WX3022,WX3008,WX2994
	,WX2980,WX2966,WX2952,WX2938,WX2924,WX2910,WX2896,WX2882
	,WX2868,WX2854,WX2840,WX2826,WX2812,WX2798,WX2784,WX2770
	,WX2756,WX2742,WX2728,WX2714,WX2700,WX2686,WX2672,WX2658
	,WX2644,WX2630,WX1771,WX1757,WX1743,WX1729,WX1715,WX1701
	,WX1687,WX1673,WX1659,WX1645,WX1631,WX1617,WX1603,WX1589
	,WX1575,WX1561,WX1547,WX1533,WX1519,WX1505,WX1491,WX1477
	,WX1463,WX1449,WX1435,WX1421,WX1407,WX1393,WX1379,WX1365
	,WX1351,WX1337,WX478,WX464,WX450,WX436,WX422,WX408
	,WX394,WX380,WX366,WX352,WX338,WX324,WX310,WX296
	,WX282,WX268,WX254,WX240,WX226,WX212,WX198,WX184
	,WX170,WX156,WX142,WX128,WX114,WX100,WX86,WX72
	,WX58,WX44,WX40,WX54,WX68,WX82,WX96,WX110
	,WX124,WX138,WX152,WX166,WX180,WX194,WX208,WX222
	,WX236,WX250,WX264,WX278,WX292,WX306,WX320,WX334
	,WX348,WX362,WX376,WX390,WX404,WX418,WX432,WX446
	,WX460,WX474,WX1333,WX1347,WX1361,WX1375,WX1389,WX1403
	,WX1417,WX1431,WX1445,WX1459,WX1473,WX1487,WX1501,WX1515
	,WX1529,WX1543,WX1557,WX1571,WX1585,WX1599,WX1613,WX1627
	,WX1641,WX1655,WX1669,WX1683,WX1697,WX1711,WX1725,WX1739
	,WX1753,WX1767,WX2626,WX2640,WX2654,WX2668,WX2682,WX2696
	,WX2710,WX2724,WX2738,WX2752,WX2766,WX2780,WX2794,WX2808
	,WX2822,WX2836,WX2850,WX2864,WX2878,WX2892,WX2906,WX2920
	,WX2934,WX2948,WX2962,WX2976,WX2990,WX3004,WX3018,WX3032
	,WX3046,WX3060,WX3919,WX3933,WX3947,WX3961,WX3975,WX3989
	,WX4003,WX4017,WX4031,WX4045,WX4059,WX4073,WX4087,WX4101
	,WX4115,WX4129,WX4143,WX4157,WX4171,WX4185,WX4199,WX4213
	,WX4227,WX4241,WX4255,WX4269,WX4283,WX4297,WX4311,WX4325
	,WX4339,WX4353,WX5212,WX5226,WX5240,WX5254,WX5268,WX5282
	,WX5296,WX5310,WX5324,WX5338,WX5352,WX5366,WX5380,WX5394
	,WX5408,WX5422,WX5436,WX5450,WX5464,WX5478,WX5492,WX5506
	,WX5520,WX5534,WX5548,WX5562,WX5576,WX5590,WX5604,WX5618
	,WX5632,WX5646,WX6505,WX6519,WX6533,WX6547,WX6561,WX6575
	,WX6589,WX6603,WX6617,WX6631,WX6645,WX6659,WX6673,WX6687
	,WX6701,WX6715,WX6729,WX6743,WX6757,WX6771,WX6785,WX6799
	,WX6813,WX6827,WX6841,WX6855,WX6869,WX6883,WX6897,WX6911
	,WX6925,WX6939,WX7798,WX7812,WX7826,WX7840,WX7854,WX7868
	,WX7882,WX7896,WX7910,WX7924,WX7938,WX7952,WX7966,WX7980
	,WX7994,WX8008,WX8022,WX8036,WX8050,WX8064,WX8078,WX8092
	,WX8106,WX8120,WX8134,WX8148,WX8162,WX8176,WX8190,WX8204
	,WX8218,WX8232,WX9091,WX9105,WX9119,WX9133,WX9147,WX9161
	,WX9175,WX9189,WX9203,WX9217,WX9231,WX9245,WX9259,WX9273
	,WX9287,WX9301,WX9315,WX9329,WX9343,WX9357,WX9371,WX9385
	,WX9399,WX9413,WX9427,WX9441,WX9455,WX9469,WX9483,WX9497
	,WX9511,WX9525,WX10824,WX10810,WX10796,WX10782,WX10768,WX10754
	,WX10740,WX10726,WX10712,WX10698,WX10684,WX10670,WX10656,WX10642
	,WX10628,WX10614,WX10600,WX10586,WX10572,WX10558,WX10544,WX10530
	,WX10516,WX10502,WX10488,WX10474,WX10460,WX10446,WX10432,WX10418
	,WX10404,WX10390,WX9531,WX9517,WX9503,WX9489,WX9475,WX9461
	,WX9447,WX9433,WX9419,WX9405,WX9391,WX9377,WX9363,WX9349
	,WX9335,WX9321,WX9307,WX9293,WX9279,WX9265,WX9251,WX9237
	,WX9223,WX9209,WX9195,WX9181,WX9167,WX9153,WX9139,WX9125
	,WX9111,WX9097,WX8238,WX8224,WX8210,WX8196,WX8182,WX8168
	,WX8154,WX8140,WX8126,WX8112,WX8098,WX8084,WX8070,WX8056
	,WX8042,WX8028,WX8014,WX8000,WX7986,WX7972,WX7958,WX7944
	,WX7930,WX7916,WX7902,WX7888,WX7874,WX7860,WX7846,WX7832
	,WX7818,WX7804,WX6945,WX6931,WX6917,WX6903,WX6889,WX6875
	,WX6861,WX6847,WX6833,WX6819,WX6805,WX6791,WX6777,WX6763
	,WX6749,WX6735,WX6721,WX6707,WX6693,WX6679,WX6665,WX6651
	,WX6637,WX6623,WX6609,WX6595,WX6581,WX6567,WX6553,WX6539
	,WX6525,WX6511,WX5652,WX5638,WX5624,WX5610,WX5596,WX5582
	,WX5568,WX5554,WX5540,WX5526,WX5512,WX5498,WX5484,WX5470
	,WX5456,WX5442,WX5428,WX5414,WX5400,WX5386,WX5372,WX5358
	,WX5344,WX5330,WX5316,WX5302,WX5288,WX5274,WX5260,WX5246
	,WX5232,WX5218,WX4359,WX4345,WX4331,WX4317,WX4303,WX4289
	,WX4275,WX4261,WX4247,WX4233,WX4219,WX4205,WX4191,WX4177
	,WX4163,WX4149,WX4135,WX4121,WX4107,WX4093,WX4079,WX4065
	,WX4051,WX4037,WX4023,WX4009,WX3995,WX3981,WX3967,WX3953
	,WX3939,WX3925,WX3066,WX3052,WX3038,WX3024,WX3010,WX2996
	,WX2982,WX2968,WX2954,WX2940,WX2926,WX2912,WX2898,WX2884
	,WX2870,WX2856,WX2842,WX2828,WX2814,WX2800,WX2786,WX2772
	,WX2758,WX2744,WX2730,WX2716,WX2702,WX2688,WX2674,WX2660
	,WX2646,WX2632,WX1773,WX1759,WX1745,WX1731,WX1717,WX1703
	,WX1689,WX1675,WX1661,WX1647,WX1633,WX1619,WX1605,WX1591
	,WX1577,WX1563,WX1549,WX1535,WX1521,WX1507,WX1493,WX1479
	,WX1465,WX1451,WX1437,WX1423,WX1409,WX1395,WX1381,WX1367
	,WX1353,WX1339,WX480,WX466,WX452,WX438,WX424,WX410
	,WX396,WX382,WX368,WX354,WX340,WX326,WX312,WX298
	,WX284,WX270,WX256,WX242,WX228,WX214,WX200,WX186
	,WX172,WX158,WX144,WX130,WX116,WX102,WX88,WX74
	,WX60,WX46,WX9093,WX9107,WX9121,WX9135,WX9149,WX9163
	,WX9177,WX9191,WX9205,WX9219,WX9233,WX9247,WX9261,WX9275
	,WX9289,WX9303,WX9317,WX9331,WX9345,WX9359,WX9373,WX9387
	,WX9401,WX9415,WX9429,WX9443,WX9457,WX9471,WX9485,WX9499
	,WX9513,WX9527,WX7800,WX7814,WX7828,WX7842,WX7856,WX7870
	,WX7884,WX7898,WX7912,WX7926,WX7940,WX7954,WX7968,WX7982
	,WX7996,WX8010,WX8024,WX8038,WX8052,WX8066,WX8080,WX8094
	,WX8108,WX8122,WX8136,WX8150,WX8164,WX8178,WX8192,WX8206
	,WX8220,WX8234,WX6507,WX6521,WX6535,WX6549,WX6563,WX6577
	,WX6591,WX6605,WX6619,WX6633,WX6647,WX6661,WX6675,WX6689
	,WX6703,WX6717,WX6731,WX6745,WX6759,WX6773,WX6787,WX6801
	,WX6815,WX6829,WX6843,WX6857,WX6871,WX6885,WX6899,WX6913
	,WX6927,WX6941,WX5214,WX5228,WX5242,WX5256,WX5270,WX5284
	,WX5298,WX5312,WX5326,WX5340,WX5354,WX5368,WX5382,WX5396
	,WX5410,WX5424,WX5438,WX5452,WX5466,WX5480,WX5494,WX5508
	,WX5522,WX5536,WX5550,WX5564,WX5578,WX5592,WX5606,WX5620
	,WX5634,WX5648,WX3921,WX3935,WX3949,WX3963,WX3977,WX3991
	,WX4005,WX4019,WX4033,WX4047,WX4061,WX4075,WX4089,WX4103
	,WX4117,WX4131,WX4145,WX4159,WX4173,WX4187,WX4201,WX4215
	,WX4229,WX4243,WX4257,WX4271,WX4285,WX4299,WX4313,WX4327
	,WX4341,WX4355,WX2628,WX2642,WX2656,WX2670,WX2684,WX2698
	,WX2712,WX2726,WX2740,WX2754,WX2768,WX2782,WX2796,WX2810
	,WX2824,WX2838,WX2852,WX2866,WX2880,WX2894,WX2908,WX2922
	,WX2936,WX2950,WX2964,WX2978,WX2992,WX3006,WX3020,WX3034
	,WX3048,WX3062,WX1335,WX1349,WX1363,WX1377,WX1391,WX1405
	,WX1419,WX1433,WX1447,WX1461,WX1475,WX1489,WX1503,WX1517
	,WX1531,WX1545,WX1559,WX1573,WX1587,WX1601,WX1615,WX1629
	,WX1643,WX1657,WX1671,WX1685,WX1699,WX1713,WX1727,WX1741
	,WX1755,WX1769,WX42,WX56,WX70,WX84,WX98,WX112
	,WX126,WX140,WX154,WX168,WX182,WX196,WX210,WX224
	,WX238,WX252,WX266,WX280,WX294,WX308,WX322,WX336
	,WX350,WX364,WX378,WX392,WX406,WX420,WX434,WX448
	,WX462,WX476,WX10813,WX10799,WX10785,WX10771,WX10757,WX10743
	,WX10729,WX10715,WX10701,WX10687,WX10673,WX10659,WX10645,WX10631
	,WX10617,WX10603,WX10589,WX10575,WX10561,WX10547,WX10533,WX10519
	,WX10505,WX10491,WX10477,WX10463,WX10449,WX10435,WX10421,WX10407
	,WX10393,WX10379,WX9520,WX9506,WX9492,WX9478,WX9464,WX9450
	,WX9436,WX9422,WX9408,WX9394,WX9380,WX9366,WX9352,WX9338
	,WX9324,WX9310,WX9296,WX9282,WX9268,WX9254,WX9240,WX9226
	,WX9212,WX9198,WX9184,WX9170,WX9156,WX9142,WX9128,WX9114
	,WX9100,WX9086,WX8227,WX8213,WX8199,WX8185,WX8171,WX8157
	,WX8143,WX8129,WX8115,WX8101,WX8087,WX8073,WX8059,WX8045
	,WX8031,WX8017,WX8003,WX7989,WX7975,WX7961,WX7947,WX7933
	,WX7919,WX7905,WX7891,WX7877,WX7863,WX7849,WX7835,WX7821
	,WX7807,WX7793,WX6934,WX6920,WX6906,WX6892,WX6878,WX6864
	,WX6850,WX6836,WX6822,WX6808,WX6794,WX6780,WX6766,WX6752
	,WX6738,WX6724,WX6710,WX6696,WX6682,WX6668,WX6654,WX6640
	,WX6626,WX6612,WX6598,WX6584,WX6570,WX6556,WX6542,WX6528
	,WX6514,WX6500,WX5641,WX5627,WX5613,WX5599,WX5585,WX5571
	,WX5557,WX5543,WX5529,WX5515,WX5501,WX5487,WX5473,WX5459
	,WX5445,WX5431,WX5417,WX5403,WX5389,WX5375,WX5361,WX5347
	,WX5333,WX5319,WX5305,WX5291,WX5277,WX5263,WX5249,WX5235
	,WX5221,WX5207,WX4348,WX4334,WX4320,WX4306,WX4292,WX4278
	,WX4264,WX4250,WX4236,WX4222,WX4208,WX4194,WX4180,WX4166
	,WX4152,WX4138,WX4124,WX4110,WX4096,WX4082,WX4068,WX4054
	,WX4040,WX4026,WX4012,WX3998,WX3984,WX3970,WX3956,WX3942
	,WX3928,WX3914,WX3055,WX3041,WX3027,WX3013,WX2999,WX2985
	,WX2971,WX2957,WX2943,WX2929,WX2915,WX2901,WX2887,WX2873
	,WX2859,WX2845,WX2831,WX2817,WX2803,WX2789,WX2775,WX2761
	,WX2747,WX2733,WX2719,WX2705,WX2691,WX2677,WX2663,WX2649
	,WX2635,WX2621,WX1762,WX1748,WX1734,WX1720,WX1706,WX1692
	,WX1678,WX1664,WX1650,WX1636,WX1622,WX1608,WX1594,WX1580
	,WX1566,WX1552,WX1538,WX1524,WX1510,WX1496,WX1482,WX1468
	,WX1454,WX1440,WX1426,WX1412,WX1398,WX1384,WX1370,WX1356
	,WX1342,WX1328,WX469,WX455,WX441,WX427,WX413,WX399
	,WX385,WX371,WX357,WX343,WX329,WX315,WX301,WX287
	,WX273,WX259,WX245,WX231,WX217,WX203,WX189,WX175
	,WX161,WX147,WX133,WX119,WX105,WX91,WX77,WX63
	,WX49,WX35,WX9521,WX9507,WX9493,WX9479,WX9465,WX9451
	,WX9437,WX9423,WX9409,WX9395,WX9381,WX9367,WX9353,WX9339
	,WX9325,WX9311,WX9297,WX9283,WX9269,WX9255,WX9241,WX9227
	,WX9213,WX9199,WX9185,WX9171,WX9157,WX9143,WX9129,WX9115
	,WX9101,WX9087,WX8228,WX8214,WX8200,WX8186,WX8172,WX8158
	,WX8144,WX8130,WX8116,WX8102,WX8088,WX8074,WX8060,WX8046
	,WX8032,WX8018,WX8004,WX7990,WX7976,WX7962,WX7948,WX7934
	,WX7920,WX7906,WX7892,WX7878,WX7864,WX7850,WX7836,WX7822
	,WX7808,WX7794,WX6935,WX6921,WX6907,WX6893,WX6879,WX6865
	,WX6851,WX6837,WX6823,WX6809,WX6795,WX6781,WX6767,WX6753
	,WX6739,WX6725,WX6711,WX6697,WX6683,WX6669,WX6655,WX6641
	,WX6627,WX6613,WX6599,WX6585,WX6571,WX6557,WX6543,WX6529
	,WX6515,WX6501,WX5642,WX5628,WX5614,WX5600,WX5586,WX5572
	,WX5558,WX5544,WX5530,WX5516,WX5502,WX5488,WX5474,WX5460
	,WX5446,WX5432,WX5418,WX5404,WX5390,WX5376,WX5362,WX5348
	,WX5334,WX5320,WX5306,WX5292,WX5278,WX5264,WX5250,WX5236
	,WX5222,WX5208,WX4349,WX4335,WX4321,WX4307,WX4293,WX4279
	,WX4265,WX4251,WX4237,WX4223,WX4209,WX4195,WX4181,WX4167
	,WX4153,WX4139,WX4125,WX4111,WX4097,WX4083,WX4069,WX4055
	,WX4041,WX4027,WX4013,WX3999,WX3985,WX3971,WX3957,WX3943
	,WX3929,WX3915,WX3056,WX3042,WX3028,WX3014,WX3000,WX2986
	,WX2972,WX2958,WX2944,WX2930,WX2916,WX2902,WX2888,WX2874
	,WX2860,WX2846,WX2832,WX2818,WX2804,WX2790,WX2776,WX2762
	,WX2748,WX2734,WX2720,WX2706,WX2692,WX2678,WX2664,WX2650
	,WX2636,WX2622,WX1763,WX1749,WX1735,WX1721,WX1707,WX1693
	,WX1679,WX1665,WX1651,WX1637,WX1623,WX1609,WX1595,WX1581
	,WX1567,WX1553,WX1539,WX1525,WX1511,WX1497,WX1483,WX1469
	,WX1455,WX1441,WX1427,WX1413,WX1399,WX1385,WX1371,WX1357
	,WX1343,WX1329,WX470,WX456,WX442,WX428,WX414,WX400
	,WX386,WX372,WX358,WX344,WX330,WX316,WX302,WX288
	,WX274,WX260,WX246,WX232,WX218,WX204,WX190,WX176
	,WX162,WX148,WX134,WX120,WX106,WX92,WX78,WX64
	,WX50,WX36,WX38,WX52,WX66,WX80,WX94,WX108
	,WX122,WX136,WX150,WX164,WX178,WX192,WX206,WX220
	,WX234,WX248,WX262,WX276,WX290,WX304,WX318,WX332
	,WX346,WX360,WX374,WX388,WX402,WX416,WX430,WX444
	,WX458,WX472,WX1331,WX1345,WX1359,WX1373,WX1387,WX1401
	,WX1415,WX1429,WX1443,WX1457,WX1471,WX1485,WX1499,WX1513
	,WX1527,WX1541,WX1555,WX1569,WX1583,WX1597,WX1611,WX1625
	,WX1639,WX1653,WX1667,WX1681,WX1695,WX1709,WX1723,WX1737
	,WX1751,WX1765,WX2624,WX2638,WX2652,WX2666,WX2680,WX2694
	,WX2708,WX2722,WX2736,WX2750,WX2764,WX2778,WX2792,WX2806
	,WX2820,WX2834,WX2848,WX2862,WX2876,WX2890,WX2904,WX2918
	,WX2932,WX2946,WX2960,WX2974,WX2988,WX3002,WX3016,WX3030
	,WX3044,WX3058,WX3917,WX3931,WX3945,WX3959,WX3973,WX3987
	,WX4001,WX4015,WX4029,WX4043,WX4057,WX4071,WX4085,WX4099
	,WX4113,WX4127,WX4141,WX4155,WX4169,WX4183,WX4197,WX4211
	,WX4225,WX4239,WX4253,WX4267,WX4281,WX4295,WX4309,WX4323
	,WX4337,WX4351,WX5210,WX5224,WX5238,WX5252,WX5266,WX5280
	,WX5294,WX5308,WX5322,WX5336,WX5350,WX5364,WX5378,WX5392
	,WX5406,WX5420,WX5434,WX5448,WX5462,WX5476,WX5490,WX5504
	,WX5518,WX5532,WX5546,WX5560,WX5574,WX5588,WX5602,WX5616
	,WX5630,WX5644,WX6503,WX6517,WX6531,WX6545,WX6559,WX6573
	,WX6587,WX6601,WX6615,WX6629,WX6643,WX6657,WX6671,WX6685
	,WX6699,WX6713,WX6727,WX6741,WX6755,WX6769,WX6783,WX6797
	,WX6811,WX6825,WX6839,WX6853,WX6867,WX6881,WX6895,WX6909
	,WX6923,WX6937,WX7796,WX7810,WX7824,WX7838,WX7852,WX7866
	,WX7880,WX7894,WX7908,WX7922,WX7936,WX7950,WX7964,WX7978
	,WX7992,WX8006,WX8020,WX8034,WX8048,WX8062,WX8076,WX8090
	,WX8104,WX8118,WX8132,WX8146,WX8160,WX8174,WX8188,WX8202
	,WX8216,WX8230,WX9089,WX9103,WX9117,WX9131,WX9145,WX9159
	,WX9173,WX9187,WX9201,WX9215,WX9229,WX9243,WX9257,WX9271
	,WX9285,WX9299,WX9313,WX9327,WX9341,WX9355,WX9369,WX9383
	,WX9397,WX9411,WX9425,WX9439,WX9453,WX9467,WX9481,WX9495
	,WX9509,WX9523,WX10382,WX10396,WX10410,WX10424,WX10438,WX10452
	,WX10466,WX10480,WX10494,WX10508,WX10522,WX10536,WX10550,WX10564
	,WX10578,WX10592,WX10606,WX10620,WX10634,WX10648,WX10662,WX10676
	,WX10690,WX10704,WX10718,WX10732,WX10746,WX10760,WX10774,WX10788
	,WX10802,WX10816,WX10825,WX10811,WX10797,WX10783,WX10769,WX10755
	,WX10741,WX10727,WX10713,WX10699,WX10685,WX10671,WX10657,WX10643
	,WX10629,WX10615,WX10601,WX10587,WX10573,WX10559,WX10545,WX10531
	,WX10517,WX10503,WX10489,WX10475,WX10461,WX10447,WX10433,WX10419
	,WX10405,WX10391,WX9532,WX9518,WX9504,WX9490,WX9476,WX9462
	,WX9448,WX9434,WX9420,WX9406,WX9392,WX9378,WX9364,WX9350
	,WX9336,WX9322,WX9308,WX9294,WX9280,WX9266,WX9252,WX9238
	,WX9224,WX9210,WX9196,WX9182,WX9168,WX9154,WX9140,WX9126
	,WX9112,WX9098,WX8239,WX8225,WX8211,WX8197,WX8183,WX8169
	,WX8155,WX8141,WX8127,WX8113,WX8099,WX8085,WX8071,WX8057
	,WX8043,WX8029,WX8015,WX8001,WX7987,WX7973,WX7959,WX7945
	,WX7931,WX7917,WX7903,WX7889,WX7875,WX7861,WX7847,WX7833
	,WX7819,WX7805,WX6946,WX6932,WX6918,WX6904,WX6890,WX6876
	,WX6862,WX6848,WX6834,WX6820,WX6806,WX6792,WX6778,WX6764
	,WX6750,WX6736,WX6722,WX6708,WX6694,WX6680,WX6666,WX6652
	,WX6638,WX6624,WX6610,WX6596,WX6582,WX6568,WX6554,WX6540
	,WX6526,WX6512,WX5653,WX5639,WX5625,WX5611,WX5597,WX5583
	,WX5569,WX5555,WX5541,WX5527,WX5513,WX5499,WX5485,WX5471
	,WX5457,WX5443,WX5429,WX5415,WX5401,WX5387,WX5373,WX5359
	,WX5345,WX5331,WX5317,WX5303,WX5289,WX5275,WX5261,WX5247
	,WX5233,WX5219,WX4360,WX4346,WX4332,WX4318,WX4304,WX4290
	,WX4276,WX4262,WX4248,WX4234,WX4220,WX4206,WX4192,WX4178
	,WX4164,WX4150,WX4136,WX4122,WX4108,WX4094,WX4080,WX4066
	,WX4052,WX4038,WX4024,WX4010,WX3996,WX3982,WX3968,WX3954
	,WX3940,WX3926,WX3067,WX3053,WX3039,WX3025,WX3011,WX2997
	,WX2983,WX2969,WX2955,WX2941,WX2927,WX2913,WX2899,WX2885
	,WX2871,WX2857,WX2843,WX2829,WX2815,WX2801,WX2787,WX2773
	,WX2759,WX2745,WX2731,WX2717,WX2703,WX2689,WX2675,WX2661
	,WX2647,WX2633,WX1774,WX1760,WX1746,WX1732,WX1718,WX1704
	,WX1690,WX1676,WX1662,WX1648,WX1634,WX1620,WX1606,WX1592
	,WX1578,WX1564,WX1550,WX1536,WX1522,WX1508,WX1494,WX1480
	,WX1466,WX1452,WX1438,WX1424,WX1410,WX1396,WX1382,WX1368
	,WX1354,WX1340,WX481,WX467,WX453,WX439,WX425,WX411
	,WX397,WX383,WX369,WX355,WX341,WX327,WX313,WX299
	,WX285,WX271,WX257,WX243,WX229,WX215,WX201,WX187
	,WX173,WX159,WX145,WX131,WX117,WX103,WX89,WX75
	,WX61,WX47,WX48,WX62,WX76,WX90,WX104,WX118
	,WX132,WX146,WX160,WX174,WX188,WX202,WX216,WX230
	,WX244,WX258,WX272,WX286,WX300,WX314,WX328,WX342
	,WX356,WX370,WX384,WX398,WX412,WX426,WX440,WX454
	,WX468,WX482,WX1341,WX1355,WX1369,WX1383,WX1397,WX1411
	,WX1425,WX1439,WX1453,WX1467,WX1481,WX1495,WX1509,WX1523
	,WX1537,WX1551,WX1565,WX1579,WX1593,WX1607,WX1621,WX1635
	,WX1649,WX1663,WX1677,WX1691,WX1705,WX1719,WX1733,WX1747
	,WX1761,WX1775,WX2634,WX2648,WX2662,WX2676,WX2690,WX2704
	,WX2718,WX2732,WX2746,WX2760,WX2774,WX2788,WX2802,WX2816
	,WX2830,WX2844,WX2858,WX2872,WX2886,WX2900,WX2914,WX2928
	,WX2942,WX2956,WX2970,WX2984,WX2998,WX3012,WX3026,WX3040
	,WX3054,WX3068,WX3927,WX3941,WX3955,WX3969,WX3983,WX3997
	,WX4011,WX4025,WX4039,WX4053,WX4067,WX4081,WX4095,WX4109
	,WX4123,WX4137,WX4151,WX4165,WX4179,WX4193,WX4207,WX4221
	,WX4235,WX4249,WX4263,WX4277,WX4291,WX4305,WX4319,WX4333
	,WX4347,WX4361,WX5220,WX5234,WX5248,WX5262,WX5276,WX5290
	,WX5304,WX5318,WX5332,WX5346,WX5360,WX5374,WX5388,WX5402
	,WX5416,WX5430,WX5444,WX5458,WX5472,WX5486,WX5500,WX5514
	,WX5528,WX5542,WX5556,WX5570,WX5584,WX5598,WX5612,WX5626
	,WX5640,WX5654,WX6513,WX6527,WX6541,WX6555,WX6569,WX6583
	,WX6597,WX6611,WX6625,WX6639,WX6653,WX6667,WX6681,WX6695
	,WX6709,WX6723,WX6737,WX6751,WX6765,WX6779,WX6793,WX6807
	,WX6821,WX6835,WX6849,WX6863,WX6877,WX6891,WX6905,WX6919
	,WX6933,WX6947,WX7806,WX7820,WX7834,WX7848,WX7862,WX7876
	,WX7890,WX7904,WX7918,WX7932,WX7946,WX7960,WX7974,WX7988
	,WX8002,WX8016,WX8030,WX8044,WX8058,WX8072,WX8086,WX8100
	,WX8114,WX8128,WX8142,WX8156,WX8170,WX8184,WX8198,WX8212
	,WX8226,WX8240,WX9099,WX9113,WX9127,WX9141,WX9155,WX9169
	,WX9183,WX9197,WX9211,WX9225,WX9239,WX9253,WX9267,WX9281
	,WX9295,WX9309,WX9323,WX9337,WX9351,WX9365,WX9379,WX9393
	,WX9407,WX9421,WX9435,WX9449,WX9463,WX9477,WX9491,WX9505
	,WX9519,WX9533,WX10392,WX10406,WX10420,WX10434,WX10448,WX10462
	,WX10476,WX10490,WX10504,WX10518,WX10532,WX10546,WX10560,WX10574
	,WX10588,WX10602,WX10616,WX10630,WX10644,WX10658,WX10672,WX10686
	,WX10700,WX10714,WX10728,WX10742,WX10756,WX10770,WX10784,WX10798
	,WX10812,WX10826,WX11050,WX11048,WX11046,WX11044,WX11042,WX11040
	,WX11038,WX11036,WX11034,WX11032,WX11030,WX11028,WX11026,WX11024
	,WX11022,WX11020,WX11018,WX11016,WX11014,WX11012,WX11010,WX11008
	,WX11006,WX11004,WX11002,WX11000,WX10998,WX10996,WX10994,WX10992
	,WX10990,WX10988,WX9757,WX9755,WX9753,WX9751,WX9749,WX9747
	,WX9745,WX9743,WX9741,WX9739,WX9737,WX9735,WX9733,WX9731
	,WX9729,WX9727,WX9725,WX9723,WX9721,WX9719,WX9717,WX9715
	,WX9713,WX9711,WX9709,WX9707,WX9705,WX9703,WX9701,WX9699
	,WX9697,WX9695,WX8464,WX8462,WX8460,WX8458,WX8456,WX8454
	,WX8452,WX8450,WX8448,WX8446,WX8444,WX8442,WX8440,WX8438
	,WX8436,WX8434,WX8432,WX8430,WX8428,WX8426,WX8424,WX8422
	,WX8420,WX8418,WX8416,WX8414,WX8412,WX8410,WX8408,WX8406
	,WX8404,WX8402,WX7171,WX7169,WX7167,WX7165,WX7163,WX7161
	,WX7159,WX7157,WX7155,WX7153,WX7151,WX7149,WX7147,WX7145
	,WX7143,WX7141,WX7139,WX7137,WX7135,WX7133,WX7131,WX7129
	,WX7127,WX7125,WX7123,WX7121,WX7119,WX7117,WX7115,WX7113
	,WX7111,WX7109,WX5878,WX5876,WX5874,WX5872,WX5870,WX5868
	,WX5866,WX5864,WX5862,WX5860,WX5858,WX5856,WX5854,WX5852
	,WX5850,WX5848,WX5846,WX5844,WX5842,WX5840,WX5838,WX5836
	,WX5834,WX5832,WX5830,WX5828,WX5826,WX5824,WX5822,WX5820
	,WX5818,WX5816,WX4585,WX4583,WX4581,WX4579,WX4577,WX4575
	,WX4573,WX4571,WX4569,WX4567,WX4565,WX4563,WX4561,WX4559
	,WX4557,WX4555,WX4553,WX4551,WX4549,WX4547,WX4545,WX4543
	,WX4541,WX4539,WX4537,WX4535,WX4533,WX4531,WX4529,WX4527
	,WX4525,WX4523,WX3292,WX3290,WX3288,WX3286,WX3284,WX3282
	,WX3280,WX3278,WX3276,WX3274,WX3272,WX3270,WX3268,WX3266
	,WX3264,WX3262,WX3260,WX3258,WX3256,WX3254,WX3252,WX3250
	,WX3248,WX3246,WX3244,WX3242,WX3240,WX3238,WX3236,WX3234
	,WX3232,WX3230,WX1999,WX1997,WX1995,WX1993,WX1991,WX1989
	,WX1987,WX1985,WX1983,WX1981,WX1979,WX1977,WX1975,WX1973
	,WX1971,WX1969,WX1967,WX1965,WX1963,WX1961,WX1959,WX1957
	,WX1955,WX1953,WX1951,WX1949,WX1947,WX1945,WX1943,WX1941
	,WX1939,WX1937,WX706,WX704,WX702,WX700,WX698,WX696
	,WX694,WX692,WX690,WX688,WX686,WX684,WX682,WX680
	,WX678,WX676,WX674,WX672,WX670,WX668,WX666,WX664
	,WX662,WX660,WX658,WX656,WX654,WX652,WX650,WX648
	,WX646,WX644;

	dff 	XG1 	(CRC_OUT_9_0,WX1264);
	dff 	XG2 	(CRC_OUT_9_1,WX1266);
	dff 	XG3 	(CRC_OUT_9_2,WX1268);
	dff 	XG4 	(CRC_OUT_9_3,WX1270);
	dff 	XG5 	(CRC_OUT_9_4,WX1272);
	dff 	XG6 	(CRC_OUT_9_5,WX1274);
	dff 	XG7 	(CRC_OUT_9_6,WX1276);
	dff 	XG8 	(CRC_OUT_9_7,WX1278);
	dff 	XG9 	(CRC_OUT_9_8,WX1280);
	dff 	XG10 	(CRC_OUT_9_9,WX1282);
	dff 	XG11 	(CRC_OUT_9_10,WX1284);
	dff 	XG12 	(CRC_OUT_9_11,WX1286);
	dff 	XG13 	(CRC_OUT_9_12,WX1288);
	dff 	XG14 	(CRC_OUT_9_13,WX1290);
	dff 	XG15 	(CRC_OUT_9_14,WX1292);
	dff 	XG16 	(CRC_OUT_9_15,WX1294);
	dff 	XG17 	(CRC_OUT_9_16,WX1296);
	dff 	XG18 	(CRC_OUT_9_17,WX1298);
	dff 	XG19 	(CRC_OUT_9_18,WX1300);
	dff 	XG20 	(CRC_OUT_9_19,WX1302);
	dff 	XG21 	(CRC_OUT_9_20,WX1304);
	dff 	XG22 	(CRC_OUT_9_21,WX1306);
	dff 	XG23 	(CRC_OUT_9_22,WX1308);
	dff 	XG24 	(CRC_OUT_9_23,WX1310);
	dff 	XG25 	(CRC_OUT_9_24,WX1312);
	dff 	XG26 	(CRC_OUT_9_25,WX1314);
	dff 	XG27 	(CRC_OUT_9_26,WX1316);
	dff 	XG28 	(CRC_OUT_9_27,WX1318);
	dff 	XG29 	(CRC_OUT_9_28,WX1320);
	dff 	XG30 	(CRC_OUT_9_29,WX1322);
	dff 	XG31 	(CRC_OUT_9_30,WX1324);
	dff 	XG32 	(CRC_OUT_9_31,WX1326);
	dff 	XG33 	(CRC_OUT_8_0,WX2557);
	dff 	XG34 	(CRC_OUT_8_1,WX2559);
	dff 	XG35 	(CRC_OUT_8_2,WX2561);
	dff 	XG36 	(CRC_OUT_8_3,WX2563);
	dff 	XG37 	(CRC_OUT_8_4,WX2565);
	dff 	XG38 	(CRC_OUT_8_5,WX2567);
	dff 	XG39 	(CRC_OUT_8_6,WX2569);
	dff 	XG40 	(CRC_OUT_8_7,WX2571);
	dff 	XG41 	(CRC_OUT_8_8,WX2573);
	dff 	XG42 	(CRC_OUT_8_9,WX2575);
	dff 	XG43 	(CRC_OUT_8_10,WX2577);
	dff 	XG44 	(CRC_OUT_8_11,WX2579);
	dff 	XG45 	(CRC_OUT_8_12,WX2581);
	dff 	XG46 	(CRC_OUT_8_13,WX2583);
	dff 	XG47 	(CRC_OUT_8_14,WX2585);
	dff 	XG48 	(CRC_OUT_8_15,WX2587);
	dff 	XG49 	(CRC_OUT_8_16,WX2589);
	dff 	XG50 	(CRC_OUT_8_17,WX2591);
	dff 	XG51 	(CRC_OUT_8_18,WX2593);
	dff 	XG52 	(CRC_OUT_8_19,WX2595);
	dff 	XG53 	(CRC_OUT_8_20,WX2597);
	dff 	XG54 	(CRC_OUT_8_21,WX2599);
	dff 	XG55 	(CRC_OUT_8_22,WX2601);
	dff 	XG56 	(CRC_OUT_8_23,WX2603);
	dff 	XG57 	(CRC_OUT_8_24,WX2605);
	dff 	XG58 	(CRC_OUT_8_25,WX2607);
	dff 	XG59 	(CRC_OUT_8_26,WX2609);
	dff 	XG60 	(CRC_OUT_8_27,WX2611);
	dff 	XG61 	(CRC_OUT_8_28,WX2613);
	dff 	XG62 	(CRC_OUT_8_29,WX2615);
	dff 	XG63 	(CRC_OUT_8_30,WX2617);
	dff 	XG64 	(CRC_OUT_8_31,WX2619);
	dff 	XG65 	(CRC_OUT_7_0,WX3850);
	dff 	XG66 	(CRC_OUT_7_1,WX3852);
	dff 	XG67 	(CRC_OUT_7_2,WX3854);
	dff 	XG68 	(CRC_OUT_7_3,WX3856);
	dff 	XG69 	(CRC_OUT_7_4,WX3858);
	dff 	XG70 	(CRC_OUT_7_5,WX3860);
	dff 	XG71 	(CRC_OUT_7_6,WX3862);
	dff 	XG72 	(CRC_OUT_7_7,WX3864);
	dff 	XG73 	(CRC_OUT_7_8,WX3866);
	dff 	XG74 	(CRC_OUT_7_9,WX3868);
	dff 	XG75 	(CRC_OUT_7_10,WX3870);
	dff 	XG76 	(CRC_OUT_7_11,WX3872);
	dff 	XG77 	(CRC_OUT_7_12,WX3874);
	dff 	XG78 	(CRC_OUT_7_13,WX3876);
	dff 	XG79 	(CRC_OUT_7_14,WX3878);
	dff 	XG80 	(CRC_OUT_7_15,WX3880);
	dff 	XG81 	(CRC_OUT_7_16,WX3882);
	dff 	XG82 	(CRC_OUT_7_17,WX3884);
	dff 	XG83 	(CRC_OUT_7_18,WX3886);
	dff 	XG84 	(CRC_OUT_7_19,WX3888);
	dff 	XG85 	(CRC_OUT_7_20,WX3890);
	dff 	XG86 	(CRC_OUT_7_21,WX3892);
	dff 	XG87 	(CRC_OUT_7_22,WX3894);
	dff 	XG88 	(CRC_OUT_7_23,WX3896);
	dff 	XG89 	(CRC_OUT_7_24,WX3898);
	dff 	XG90 	(CRC_OUT_7_25,WX3900);
	dff 	XG91 	(CRC_OUT_7_26,WX3902);
	dff 	XG92 	(CRC_OUT_7_27,WX3904);
	dff 	XG93 	(CRC_OUT_7_28,WX3906);
	dff 	XG94 	(CRC_OUT_7_29,WX3908);
	dff 	XG95 	(CRC_OUT_7_30,WX3910);
	dff 	XG96 	(CRC_OUT_7_31,WX3912);
	dff 	XG97 	(CRC_OUT_6_0,WX5143);
	dff 	XG98 	(CRC_OUT_6_1,WX5145);
	dff 	XG99 	(CRC_OUT_6_2,WX5147);
	dff 	XG100 	(CRC_OUT_6_3,WX5149);
	dff 	XG101 	(CRC_OUT_6_4,WX5151);
	dff 	XG102 	(CRC_OUT_6_5,WX5153);
	dff 	XG103 	(CRC_OUT_6_6,WX5155);
	dff 	XG104 	(CRC_OUT_6_7,WX5157);
	dff 	XG105 	(CRC_OUT_6_8,WX5159);
	dff 	XG106 	(CRC_OUT_6_9,WX5161);
	dff 	XG107 	(CRC_OUT_6_10,WX5163);
	dff 	XG108 	(CRC_OUT_6_11,WX5165);
	dff 	XG109 	(CRC_OUT_6_12,WX5167);
	dff 	XG110 	(CRC_OUT_6_13,WX5169);
	dff 	XG111 	(CRC_OUT_6_14,WX5171);
	dff 	XG112 	(CRC_OUT_6_15,WX5173);
	dff 	XG113 	(CRC_OUT_6_16,WX5175);
	dff 	XG114 	(CRC_OUT_6_17,WX5177);
	dff 	XG115 	(CRC_OUT_6_18,WX5179);
	dff 	XG116 	(CRC_OUT_6_19,WX5181);
	dff 	XG117 	(CRC_OUT_6_20,WX5183);
	dff 	XG118 	(CRC_OUT_6_21,WX5185);
	dff 	XG119 	(CRC_OUT_6_22,WX5187);
	dff 	XG120 	(CRC_OUT_6_23,WX5189);
	dff 	XG121 	(CRC_OUT_6_24,WX5191);
	dff 	XG122 	(CRC_OUT_6_25,WX5193);
	dff 	XG123 	(CRC_OUT_6_26,WX5195);
	dff 	XG124 	(CRC_OUT_6_27,WX5197);
	dff 	XG125 	(CRC_OUT_6_28,WX5199);
	dff 	XG126 	(CRC_OUT_6_29,WX5201);
	dff 	XG127 	(CRC_OUT_6_30,WX5203);
	dff 	XG128 	(CRC_OUT_6_31,WX5205);
	dff 	XG129 	(CRC_OUT_5_0,WX6436);
	dff 	XG130 	(CRC_OUT_5_1,WX6438);
	dff 	XG131 	(CRC_OUT_5_2,WX6440);
	dff 	XG132 	(CRC_OUT_5_3,WX6442);
	dff 	XG133 	(CRC_OUT_5_4,WX6444);
	dff 	XG134 	(CRC_OUT_5_5,WX6446);
	dff 	XG135 	(CRC_OUT_5_6,WX6448);
	dff 	XG136 	(CRC_OUT_5_7,WX6450);
	dff 	XG137 	(CRC_OUT_5_8,WX6452);
	dff 	XG138 	(CRC_OUT_5_9,WX6454);
	dff 	XG139 	(CRC_OUT_5_10,WX6456);
	dff 	XG140 	(CRC_OUT_5_11,WX6458);
	dff 	XG141 	(CRC_OUT_5_12,WX6460);
	dff 	XG142 	(CRC_OUT_5_13,WX6462);
	dff 	XG143 	(CRC_OUT_5_14,WX6464);
	dff 	XG144 	(CRC_OUT_5_15,WX6466);
	dff 	XG145 	(CRC_OUT_5_16,WX6468);
	dff 	XG146 	(CRC_OUT_5_17,WX6470);
	dff 	XG147 	(CRC_OUT_5_18,WX6472);
	dff 	XG148 	(CRC_OUT_5_19,WX6474);
	dff 	XG149 	(CRC_OUT_5_20,WX6476);
	dff 	XG150 	(CRC_OUT_5_21,WX6478);
	dff 	XG151 	(CRC_OUT_5_22,WX6480);
	dff 	XG152 	(CRC_OUT_5_23,WX6482);
	dff 	XG153 	(CRC_OUT_5_24,WX6484);
	dff 	XG154 	(CRC_OUT_5_25,WX6486);
	dff 	XG155 	(CRC_OUT_5_26,WX6488);
	dff 	XG156 	(CRC_OUT_5_27,WX6490);
	dff 	XG157 	(CRC_OUT_5_28,WX6492);
	dff 	XG158 	(CRC_OUT_5_29,WX6494);
	dff 	XG159 	(CRC_OUT_5_30,WX6496);
	dff 	XG160 	(CRC_OUT_5_31,WX6498);
	dff 	XG161 	(CRC_OUT_4_0,WX7729);
	dff 	XG162 	(CRC_OUT_4_1,WX7731);
	dff 	XG163 	(CRC_OUT_4_2,WX7733);
	dff 	XG164 	(CRC_OUT_4_3,WX7735);
	dff 	XG165 	(CRC_OUT_4_4,WX7737);
	dff 	XG166 	(CRC_OUT_4_5,WX7739);
	dff 	XG167 	(CRC_OUT_4_6,WX7741);
	dff 	XG168 	(CRC_OUT_4_7,WX7743);
	dff 	XG169 	(CRC_OUT_4_8,WX7745);
	dff 	XG170 	(CRC_OUT_4_9,WX7747);
	dff 	XG171 	(CRC_OUT_4_10,WX7749);
	dff 	XG172 	(CRC_OUT_4_11,WX7751);
	dff 	XG173 	(CRC_OUT_4_12,WX7753);
	dff 	XG174 	(CRC_OUT_4_13,WX7755);
	dff 	XG175 	(CRC_OUT_4_14,WX7757);
	dff 	XG176 	(CRC_OUT_4_15,WX7759);
	dff 	XG177 	(CRC_OUT_4_16,WX7761);
	dff 	XG178 	(CRC_OUT_4_17,WX7763);
	dff 	XG179 	(CRC_OUT_4_18,WX7765);
	dff 	XG180 	(CRC_OUT_4_19,WX7767);
	dff 	XG181 	(CRC_OUT_4_20,WX7769);
	dff 	XG182 	(CRC_OUT_4_21,WX7771);
	dff 	XG183 	(CRC_OUT_4_22,WX7773);
	dff 	XG184 	(CRC_OUT_4_23,WX7775);
	dff 	XG185 	(CRC_OUT_4_24,WX7777);
	dff 	XG186 	(CRC_OUT_4_25,WX7779);
	dff 	XG187 	(CRC_OUT_4_26,WX7781);
	dff 	XG188 	(CRC_OUT_4_27,WX7783);
	dff 	XG189 	(CRC_OUT_4_28,WX7785);
	dff 	XG190 	(CRC_OUT_4_29,WX7787);
	dff 	XG191 	(CRC_OUT_4_30,WX7789);
	dff 	XG192 	(CRC_OUT_4_31,WX7791);
	dff 	XG193 	(CRC_OUT_3_0,WX9022);
	dff 	XG194 	(CRC_OUT_3_1,WX9024);
	dff 	XG195 	(CRC_OUT_3_2,WX9026);
	dff 	XG196 	(CRC_OUT_3_3,WX9028);
	dff 	XG197 	(CRC_OUT_3_4,WX9030);
	dff 	XG198 	(CRC_OUT_3_5,WX9032);
	dff 	XG199 	(CRC_OUT_3_6,WX9034);
	dff 	XG200 	(CRC_OUT_3_7,WX9036);
	dff 	XG201 	(CRC_OUT_3_8,WX9038);
	dff 	XG202 	(CRC_OUT_3_9,WX9040);
	dff 	XG203 	(CRC_OUT_3_10,WX9042);
	dff 	XG204 	(CRC_OUT_3_11,WX9044);
	dff 	XG205 	(CRC_OUT_3_12,WX9046);
	dff 	XG206 	(CRC_OUT_3_13,WX9048);
	dff 	XG207 	(CRC_OUT_3_14,WX9050);
	dff 	XG208 	(CRC_OUT_3_15,WX9052);
	dff 	XG209 	(CRC_OUT_3_16,WX9054);
	dff 	XG210 	(CRC_OUT_3_17,WX9056);
	dff 	XG211 	(CRC_OUT_3_18,WX9058);
	dff 	XG212 	(CRC_OUT_3_19,WX9060);
	dff 	XG213 	(CRC_OUT_3_20,WX9062);
	dff 	XG214 	(CRC_OUT_3_21,WX9064);
	dff 	XG215 	(CRC_OUT_3_22,WX9066);
	dff 	XG216 	(CRC_OUT_3_23,WX9068);
	dff 	XG217 	(CRC_OUT_3_24,WX9070);
	dff 	XG218 	(CRC_OUT_3_25,WX9072);
	dff 	XG219 	(CRC_OUT_3_26,WX9074);
	dff 	XG220 	(CRC_OUT_3_27,WX9076);
	dff 	XG221 	(CRC_OUT_3_28,WX9078);
	dff 	XG222 	(CRC_OUT_3_29,WX9080);
	dff 	XG223 	(CRC_OUT_3_30,WX9082);
	dff 	XG224 	(CRC_OUT_3_31,WX9084);
	dff 	XG225 	(CRC_OUT_2_0,WX10315);
	dff 	XG226 	(CRC_OUT_2_1,WX10317);
	dff 	XG227 	(CRC_OUT_2_2,WX10319);
	dff 	XG228 	(CRC_OUT_2_3,WX10321);
	dff 	XG229 	(CRC_OUT_2_4,WX10323);
	dff 	XG230 	(CRC_OUT_2_5,WX10325);
	dff 	XG231 	(CRC_OUT_2_6,WX10327);
	dff 	XG232 	(CRC_OUT_2_7,WX10329);
	dff 	XG233 	(CRC_OUT_2_8,WX10331);
	dff 	XG234 	(CRC_OUT_2_9,WX10333);
	dff 	XG235 	(CRC_OUT_2_10,WX10335);
	dff 	XG236 	(CRC_OUT_2_11,WX10337);
	dff 	XG237 	(CRC_OUT_2_12,WX10339);
	dff 	XG238 	(CRC_OUT_2_13,WX10341);
	dff 	XG239 	(CRC_OUT_2_14,WX10343);
	dff 	XG240 	(CRC_OUT_2_15,WX10345);
	dff 	XG241 	(CRC_OUT_2_16,WX10347);
	dff 	XG242 	(CRC_OUT_2_17,WX10349);
	dff 	XG243 	(CRC_OUT_2_18,WX10351);
	dff 	XG244 	(CRC_OUT_2_19,WX10353);
	dff 	XG245 	(CRC_OUT_2_20,WX10355);
	dff 	XG246 	(CRC_OUT_2_21,WX10357);
	dff 	XG247 	(CRC_OUT_2_22,WX10359);
	dff 	XG248 	(CRC_OUT_2_23,WX10361);
	dff 	XG249 	(CRC_OUT_2_24,WX10363);
	dff 	XG250 	(CRC_OUT_2_25,WX10365);
	dff 	XG251 	(CRC_OUT_2_26,WX10367);
	dff 	XG252 	(CRC_OUT_2_27,WX10369);
	dff 	XG253 	(CRC_OUT_2_28,WX10371);
	dff 	XG254 	(CRC_OUT_2_29,WX10373);
	dff 	XG255 	(CRC_OUT_2_30,WX10375);
	dff 	XG256 	(CRC_OUT_2_31,WX10377);
	dff 	XG257 	(CRC_OUT_1_0,WX11608);
	dff 	XG258 	(CRC_OUT_1_1,WX11610);
	dff 	XG259 	(CRC_OUT_1_2,WX11612);
	dff 	XG260 	(CRC_OUT_1_3,WX11614);
	dff 	XG261 	(CRC_OUT_1_4,WX11616);
	dff 	XG262 	(CRC_OUT_1_5,WX11618);
	dff 	XG263 	(CRC_OUT_1_6,WX11620);
	dff 	XG264 	(CRC_OUT_1_7,WX11622);
	dff 	XG265 	(CRC_OUT_1_8,WX11624);
	dff 	XG266 	(CRC_OUT_1_9,WX11626);
	dff 	XG267 	(CRC_OUT_1_10,WX11628);
	dff 	XG268 	(CRC_OUT_1_11,WX11630);
	dff 	XG269 	(CRC_OUT_1_12,WX11632);
	dff 	XG270 	(CRC_OUT_1_13,WX11634);
	dff 	XG271 	(CRC_OUT_1_14,WX11636);
	dff 	XG272 	(CRC_OUT_1_15,WX11638);
	dff 	XG273 	(CRC_OUT_1_16,WX11640);
	dff 	XG274 	(CRC_OUT_1_17,WX11642);
	dff 	XG275 	(CRC_OUT_1_18,WX11644);
	dff 	XG276 	(CRC_OUT_1_19,WX11646);
	dff 	XG277 	(CRC_OUT_1_20,WX11648);
	dff 	XG278 	(CRC_OUT_1_21,WX11650);
	dff 	XG279 	(CRC_OUT_1_22,WX11652);
	dff 	XG280 	(CRC_OUT_1_23,WX11654);
	dff 	XG281 	(CRC_OUT_1_24,WX11656);
	dff 	XG282 	(CRC_OUT_1_25,WX11658);
	dff 	XG283 	(CRC_OUT_1_26,WX11660);
	dff 	XG284 	(CRC_OUT_1_27,WX11662);
	dff 	XG285 	(CRC_OUT_1_28,WX11664);
	dff 	XG286 	(CRC_OUT_1_29,WX11666);
	dff 	XG287 	(CRC_OUT_1_30,WX11668);
	dff 	XG288 	(CRC_OUT_1_31,WX11670);
	dff 	XG289 	(WX485,WX484);
	dff 	XG290 	(WX487,WX486);
	dff 	XG291 	(WX489,WX488);
	dff 	XG292 	(WX491,WX490);
	dff 	XG293 	(WX493,WX492);
	dff 	XG294 	(WX495,WX494);
	dff 	XG295 	(WX497,WX496);
	dff 	XG296 	(WX499,WX498);
	dff 	XG297 	(WX501,WX500);
	dff 	XG298 	(WX503,WX502);
	dff 	XG299 	(WX505,WX504);
	dff 	XG300 	(WX507,WX506);
	dff 	XG301 	(WX509,WX508);
	dff 	XG302 	(WX511,WX510);
	dff 	XG303 	(WX513,WX512);
	dff 	XG304 	(WX515,WX514);
	dff 	XG305 	(WX517,WX516);
	dff 	XG306 	(WX519,WX518);
	dff 	XG307 	(WX521,WX520);
	dff 	XG308 	(WX523,WX522);
	dff 	XG309 	(WX525,WX524);
	dff 	XG310 	(WX527,WX526);
	dff 	XG311 	(WX529,WX528);
	dff 	XG312 	(WX531,WX530);
	dff 	XG313 	(WX533,WX532);
	dff 	XG314 	(WX535,WX534);
	dff 	XG315 	(WX537,WX536);
	dff 	XG316 	(WX539,WX538);
	dff 	XG317 	(WX541,WX540);
	dff 	XG318 	(WX543,WX542);
	dff 	XG319 	(WX545,WX544);
	dff 	XG320 	(WX547,WX546);
	dff 	XG321 	(WX645,WX644);
	dff 	XG322 	(WX647,WX646);
	dff 	XG323 	(WX649,WX648);
	dff 	XG324 	(WX651,WX650);
	dff 	XG325 	(WX653,WX652);
	dff 	XG326 	(WX655,WX654);
	dff 	XG327 	(WX657,WX656);
	dff 	XG328 	(WX659,WX658);
	dff 	XG329 	(WX661,WX660);
	dff 	XG330 	(WX663,WX662);
	dff 	XG331 	(WX665,WX664);
	dff 	XG332 	(WX667,WX666);
	dff 	XG333 	(WX669,WX668);
	dff 	XG334 	(WX671,WX670);
	dff 	XG335 	(WX673,WX672);
	dff 	XG336 	(WX675,WX674);
	dff 	XG337 	(WX677,WX676);
	dff 	XG338 	(WX679,WX678);
	dff 	XG339 	(WX681,WX680);
	dff 	XG340 	(WX683,WX682);
	dff 	XG341 	(WX685,WX684);
	dff 	XG342 	(WX687,WX686);
	dff 	XG343 	(WX689,WX688);
	dff 	XG344 	(WX691,WX690);
	dff 	XG345 	(WX693,WX692);
	dff 	XG346 	(WX695,WX694);
	dff 	XG347 	(WX697,WX696);
	dff 	XG348 	(WX699,WX698);
	dff 	XG349 	(WX701,WX700);
	dff 	XG350 	(WX703,WX702);
	dff 	XG351 	(WX705,WX704);
	dff 	XG352 	(WX707,WX706);
	dff 	XG353 	(WX709,WX708);
	dff 	XG354 	(WX711,WX710);
	dff 	XG355 	(WX713,WX712);
	dff 	XG356 	(WX715,WX714);
	dff 	XG357 	(WX717,WX716);
	dff 	XG358 	(WX719,WX718);
	dff 	XG359 	(WX721,WX720);
	dff 	XG360 	(WX723,WX722);
	dff 	XG361 	(WX725,WX724);
	dff 	XG362 	(WX727,WX726);
	dff 	XG363 	(WX729,WX728);
	dff 	XG364 	(WX731,WX730);
	dff 	XG365 	(WX733,WX732);
	dff 	XG366 	(WX735,WX734);
	dff 	XG367 	(WX737,WX736);
	dff 	XG368 	(WX739,WX738);
	dff 	XG369 	(WX741,WX740);
	dff 	XG370 	(WX743,WX742);
	dff 	XG371 	(WX745,WX744);
	dff 	XG372 	(WX747,WX746);
	dff 	XG373 	(WX749,WX748);
	dff 	XG374 	(WX751,WX750);
	dff 	XG375 	(WX753,WX752);
	dff 	XG376 	(WX755,WX754);
	dff 	XG377 	(WX757,WX756);
	dff 	XG378 	(WX759,WX758);
	dff 	XG379 	(WX761,WX760);
	dff 	XG380 	(WX763,WX762);
	dff 	XG381 	(WX765,WX764);
	dff 	XG382 	(WX767,WX766);
	dff 	XG383 	(WX769,WX768);
	dff 	XG384 	(WX771,WX770);
	dff 	XG385 	(WX773,WX772);
	dff 	XG386 	(WX775,WX774);
	dff 	XG387 	(WX777,WX776);
	dff 	XG388 	(WX779,WX778);
	dff 	XG389 	(WX781,WX780);
	dff 	XG390 	(WX783,WX782);
	dff 	XG391 	(WX785,WX784);
	dff 	XG392 	(WX787,WX786);
	dff 	XG393 	(WX789,WX788);
	dff 	XG394 	(WX791,WX790);
	dff 	XG395 	(WX793,WX792);
	dff 	XG396 	(WX795,WX794);
	dff 	XG397 	(WX797,WX796);
	dff 	XG398 	(WX799,WX798);
	dff 	XG399 	(WX801,WX800);
	dff 	XG400 	(WX803,WX802);
	dff 	XG401 	(WX805,WX804);
	dff 	XG402 	(WX807,WX806);
	dff 	XG403 	(WX809,WX808);
	dff 	XG404 	(WX811,WX810);
	dff 	XG405 	(WX813,WX812);
	dff 	XG406 	(WX815,WX814);
	dff 	XG407 	(WX817,WX816);
	dff 	XG408 	(WX819,WX818);
	dff 	XG409 	(WX821,WX820);
	dff 	XG410 	(WX823,WX822);
	dff 	XG411 	(WX825,WX824);
	dff 	XG412 	(WX827,WX826);
	dff 	XG413 	(WX829,WX828);
	dff 	XG414 	(WX831,WX830);
	dff 	XG415 	(WX833,WX832);
	dff 	XG416 	(WX835,WX834);
	dff 	XG417 	(WX837,WX836);
	dff 	XG418 	(WX839,WX838);
	dff 	XG419 	(WX841,WX840);
	dff 	XG420 	(WX843,WX842);
	dff 	XG421 	(WX845,WX844);
	dff 	XG422 	(WX847,WX846);
	dff 	XG423 	(WX849,WX848);
	dff 	XG424 	(WX851,WX850);
	dff 	XG425 	(WX853,WX852);
	dff 	XG426 	(WX855,WX854);
	dff 	XG427 	(WX857,WX856);
	dff 	XG428 	(WX859,WX858);
	dff 	XG429 	(WX861,WX860);
	dff 	XG430 	(WX863,WX862);
	dff 	XG431 	(WX865,WX864);
	dff 	XG432 	(WX867,WX866);
	dff 	XG433 	(WX869,WX868);
	dff 	XG434 	(WX871,WX870);
	dff 	XG435 	(WX873,WX872);
	dff 	XG436 	(WX875,WX874);
	dff 	XG437 	(WX877,WX876);
	dff 	XG438 	(WX879,WX878);
	dff 	XG439 	(WX881,WX880);
	dff 	XG440 	(WX883,WX882);
	dff 	XG441 	(WX885,WX884);
	dff 	XG442 	(WX887,WX886);
	dff 	XG443 	(WX889,WX888);
	dff 	XG444 	(WX891,WX890);
	dff 	XG445 	(WX893,WX892);
	dff 	XG446 	(WX895,WX894);
	dff 	XG447 	(WX897,WX896);
	dff 	XG448 	(WX899,WX898);
	dff 	XG449 	(WX1778,WX1777);
	dff 	XG450 	(WX1780,WX1779);
	dff 	XG451 	(WX1782,WX1781);
	dff 	XG452 	(WX1784,WX1783);
	dff 	XG453 	(WX1786,WX1785);
	dff 	XG454 	(WX1788,WX1787);
	dff 	XG455 	(WX1790,WX1789);
	dff 	XG456 	(WX1792,WX1791);
	dff 	XG457 	(WX1794,WX1793);
	dff 	XG458 	(WX1796,WX1795);
	dff 	XG459 	(WX1798,WX1797);
	dff 	XG460 	(WX1800,WX1799);
	dff 	XG461 	(WX1802,WX1801);
	dff 	XG462 	(WX1804,WX1803);
	dff 	XG463 	(WX1806,WX1805);
	dff 	XG464 	(WX1808,WX1807);
	dff 	XG465 	(WX1810,WX1809);
	dff 	XG466 	(WX1812,WX1811);
	dff 	XG467 	(WX1814,WX1813);
	dff 	XG468 	(WX1816,WX1815);
	dff 	XG469 	(WX1818,WX1817);
	dff 	XG470 	(WX1820,WX1819);
	dff 	XG471 	(WX1822,WX1821);
	dff 	XG472 	(WX1824,WX1823);
	dff 	XG473 	(WX1826,WX1825);
	dff 	XG474 	(WX1828,WX1827);
	dff 	XG475 	(WX1830,WX1829);
	dff 	XG476 	(WX1832,WX1831);
	dff 	XG477 	(WX1834,WX1833);
	dff 	XG478 	(WX1836,WX1835);
	dff 	XG479 	(WX1838,WX1837);
	dff 	XG480 	(WX1840,WX1839);
	dff 	XG481 	(WX1938,WX1937);
	dff 	XG482 	(WX1940,WX1939);
	dff 	XG483 	(WX1942,WX1941);
	dff 	XG484 	(WX1944,WX1943);
	dff 	XG485 	(WX1946,WX1945);
	dff 	XG486 	(WX1948,WX1947);
	dff 	XG487 	(WX1950,WX1949);
	dff 	XG488 	(WX1952,WX1951);
	dff 	XG489 	(WX1954,WX1953);
	dff 	XG490 	(WX1956,WX1955);
	dff 	XG491 	(WX1958,WX1957);
	dff 	XG492 	(WX1960,WX1959);
	dff 	XG493 	(WX1962,WX1961);
	dff 	XG494 	(WX1964,WX1963);
	dff 	XG495 	(WX1966,WX1965);
	dff 	XG496 	(WX1968,WX1967);
	dff 	XG497 	(WX1970,WX1969);
	dff 	XG498 	(WX1972,WX1971);
	dff 	XG499 	(WX1974,WX1973);
	dff 	XG500 	(WX1976,WX1975);
	dff 	XG501 	(WX1978,WX1977);
	dff 	XG502 	(WX1980,WX1979);
	dff 	XG503 	(WX1982,WX1981);
	dff 	XG504 	(WX1984,WX1983);
	dff 	XG505 	(WX1986,WX1985);
	dff 	XG506 	(WX1988,WX1987);
	dff 	XG507 	(WX1990,WX1989);
	dff 	XG508 	(WX1992,WX1991);
	dff 	XG509 	(WX1994,WX1993);
	dff 	XG510 	(WX1996,WX1995);
	dff 	XG511 	(WX1998,WX1997);
	dff 	XG512 	(WX2000,WX1999);
	dff 	XG513 	(WX2002,WX2001);
	dff 	XG514 	(WX2004,WX2003);
	dff 	XG515 	(WX2006,WX2005);
	dff 	XG516 	(WX2008,WX2007);
	dff 	XG517 	(WX2010,WX2009);
	dff 	XG518 	(WX2012,WX2011);
	dff 	XG519 	(WX2014,WX2013);
	dff 	XG520 	(WX2016,WX2015);
	dff 	XG521 	(WX2018,WX2017);
	dff 	XG522 	(WX2020,WX2019);
	dff 	XG523 	(WX2022,WX2021);
	dff 	XG524 	(WX2024,WX2023);
	dff 	XG525 	(WX2026,WX2025);
	dff 	XG526 	(WX2028,WX2027);
	dff 	XG527 	(WX2030,WX2029);
	dff 	XG528 	(WX2032,WX2031);
	dff 	XG529 	(WX2034,WX2033);
	dff 	XG530 	(WX2036,WX2035);
	dff 	XG531 	(WX2038,WX2037);
	dff 	XG532 	(WX2040,WX2039);
	dff 	XG533 	(WX2042,WX2041);
	dff 	XG534 	(WX2044,WX2043);
	dff 	XG535 	(WX2046,WX2045);
	dff 	XG536 	(WX2048,WX2047);
	dff 	XG537 	(WX2050,WX2049);
	dff 	XG538 	(WX2052,WX2051);
	dff 	XG539 	(WX2054,WX2053);
	dff 	XG540 	(WX2056,WX2055);
	dff 	XG541 	(WX2058,WX2057);
	dff 	XG542 	(WX2060,WX2059);
	dff 	XG543 	(WX2062,WX2061);
	dff 	XG544 	(WX2064,WX2063);
	dff 	XG545 	(WX2066,WX2065);
	dff 	XG546 	(WX2068,WX2067);
	dff 	XG547 	(WX2070,WX2069);
	dff 	XG548 	(WX2072,WX2071);
	dff 	XG549 	(WX2074,WX2073);
	dff 	XG550 	(WX2076,WX2075);
	dff 	XG551 	(WX2078,WX2077);
	dff 	XG552 	(WX2080,WX2079);
	dff 	XG553 	(WX2082,WX2081);
	dff 	XG554 	(WX2084,WX2083);
	dff 	XG555 	(WX2086,WX2085);
	dff 	XG556 	(WX2088,WX2087);
	dff 	XG557 	(WX2090,WX2089);
	dff 	XG558 	(WX2092,WX2091);
	dff 	XG559 	(WX2094,WX2093);
	dff 	XG560 	(WX2096,WX2095);
	dff 	XG561 	(WX2098,WX2097);
	dff 	XG562 	(WX2100,WX2099);
	dff 	XG563 	(WX2102,WX2101);
	dff 	XG564 	(WX2104,WX2103);
	dff 	XG565 	(WX2106,WX2105);
	dff 	XG566 	(WX2108,WX2107);
	dff 	XG567 	(WX2110,WX2109);
	dff 	XG568 	(WX2112,WX2111);
	dff 	XG569 	(WX2114,WX2113);
	dff 	XG570 	(WX2116,WX2115);
	dff 	XG571 	(WX2118,WX2117);
	dff 	XG572 	(WX2120,WX2119);
	dff 	XG573 	(WX2122,WX2121);
	dff 	XG574 	(WX2124,WX2123);
	dff 	XG575 	(WX2126,WX2125);
	dff 	XG576 	(WX2128,WX2127);
	dff 	XG577 	(WX2130,WX2129);
	dff 	XG578 	(WX2132,WX2131);
	dff 	XG579 	(WX2134,WX2133);
	dff 	XG580 	(WX2136,WX2135);
	dff 	XG581 	(WX2138,WX2137);
	dff 	XG582 	(WX2140,WX2139);
	dff 	XG583 	(WX2142,WX2141);
	dff 	XG584 	(WX2144,WX2143);
	dff 	XG585 	(WX2146,WX2145);
	dff 	XG586 	(WX2148,WX2147);
	dff 	XG587 	(WX2150,WX2149);
	dff 	XG588 	(WX2152,WX2151);
	dff 	XG589 	(WX2154,WX2153);
	dff 	XG590 	(WX2156,WX2155);
	dff 	XG591 	(WX2158,WX2157);
	dff 	XG592 	(WX2160,WX2159);
	dff 	XG593 	(WX2162,WX2161);
	dff 	XG594 	(WX2164,WX2163);
	dff 	XG595 	(WX2166,WX2165);
	dff 	XG596 	(WX2168,WX2167);
	dff 	XG597 	(WX2170,WX2169);
	dff 	XG598 	(WX2172,WX2171);
	dff 	XG599 	(WX2174,WX2173);
	dff 	XG600 	(WX2176,WX2175);
	dff 	XG601 	(WX2178,WX2177);
	dff 	XG602 	(WX2180,WX2179);
	dff 	XG603 	(WX2182,WX2181);
	dff 	XG604 	(WX2184,WX2183);
	dff 	XG605 	(WX2186,WX2185);
	dff 	XG606 	(WX2188,WX2187);
	dff 	XG607 	(WX2190,WX2189);
	dff 	XG608 	(WX2192,WX2191);
	dff 	XG609 	(WX3071,WX3070);
	dff 	XG610 	(WX3073,WX3072);
	dff 	XG611 	(WX3075,WX3074);
	dff 	XG612 	(WX3077,WX3076);
	dff 	XG613 	(WX3079,WX3078);
	dff 	XG614 	(WX3081,WX3080);
	dff 	XG615 	(WX3083,WX3082);
	dff 	XG616 	(WX3085,WX3084);
	dff 	XG617 	(WX3087,WX3086);
	dff 	XG618 	(WX3089,WX3088);
	dff 	XG619 	(WX3091,WX3090);
	dff 	XG620 	(WX3093,WX3092);
	dff 	XG621 	(WX3095,WX3094);
	dff 	XG622 	(WX3097,WX3096);
	dff 	XG623 	(WX3099,WX3098);
	dff 	XG624 	(WX3101,WX3100);
	dff 	XG625 	(WX3103,WX3102);
	dff 	XG626 	(WX3105,WX3104);
	dff 	XG627 	(WX3107,WX3106);
	dff 	XG628 	(WX3109,WX3108);
	dff 	XG629 	(WX3111,WX3110);
	dff 	XG630 	(WX3113,WX3112);
	dff 	XG631 	(WX3115,WX3114);
	dff 	XG632 	(WX3117,WX3116);
	dff 	XG633 	(WX3119,WX3118);
	dff 	XG634 	(WX3121,WX3120);
	dff 	XG635 	(WX3123,WX3122);
	dff 	XG636 	(WX3125,WX3124);
	dff 	XG637 	(WX3127,WX3126);
	dff 	XG638 	(WX3129,WX3128);
	dff 	XG639 	(WX3131,WX3130);
	dff 	XG640 	(WX3133,WX3132);
	dff 	XG641 	(WX3231,WX3230);
	dff 	XG642 	(WX3233,WX3232);
	dff 	XG643 	(WX3235,WX3234);
	dff 	XG644 	(WX3237,WX3236);
	dff 	XG645 	(WX3239,WX3238);
	dff 	XG646 	(WX3241,WX3240);
	dff 	XG647 	(WX3243,WX3242);
	dff 	XG648 	(WX3245,WX3244);
	dff 	XG649 	(WX3247,WX3246);
	dff 	XG650 	(WX3249,WX3248);
	dff 	XG651 	(WX3251,WX3250);
	dff 	XG652 	(WX3253,WX3252);
	dff 	XG653 	(WX3255,WX3254);
	dff 	XG654 	(WX3257,WX3256);
	dff 	XG655 	(WX3259,WX3258);
	dff 	XG656 	(WX3261,WX3260);
	dff 	XG657 	(WX3263,WX3262);
	dff 	XG658 	(WX3265,WX3264);
	dff 	XG659 	(WX3267,WX3266);
	dff 	XG660 	(WX3269,WX3268);
	dff 	XG661 	(WX3271,WX3270);
	dff 	XG662 	(WX3273,WX3272);
	dff 	XG663 	(WX3275,WX3274);
	dff 	XG664 	(WX3277,WX3276);
	dff 	XG665 	(WX3279,WX3278);
	dff 	XG666 	(WX3281,WX3280);
	dff 	XG667 	(WX3283,WX3282);
	dff 	XG668 	(WX3285,WX3284);
	dff 	XG669 	(WX3287,WX3286);
	dff 	XG670 	(WX3289,WX3288);
	dff 	XG671 	(WX3291,WX3290);
	dff 	XG672 	(WX3293,WX3292);
	dff 	XG673 	(WX3295,WX3294);
	dff 	XG674 	(WX3297,WX3296);
	dff 	XG675 	(WX3299,WX3298);
	dff 	XG676 	(WX3301,WX3300);
	dff 	XG677 	(WX3303,WX3302);
	dff 	XG678 	(WX3305,WX3304);
	dff 	XG679 	(WX3307,WX3306);
	dff 	XG680 	(WX3309,WX3308);
	dff 	XG681 	(WX3311,WX3310);
	dff 	XG682 	(WX3313,WX3312);
	dff 	XG683 	(WX3315,WX3314);
	dff 	XG684 	(WX3317,WX3316);
	dff 	XG685 	(WX3319,WX3318);
	dff 	XG686 	(WX3321,WX3320);
	dff 	XG687 	(WX3323,WX3322);
	dff 	XG688 	(WX3325,WX3324);
	dff 	XG689 	(WX3327,WX3326);
	dff 	XG690 	(WX3329,WX3328);
	dff 	XG691 	(WX3331,WX3330);
	dff 	XG692 	(WX3333,WX3332);
	dff 	XG693 	(WX3335,WX3334);
	dff 	XG694 	(WX3337,WX3336);
	dff 	XG695 	(WX3339,WX3338);
	dff 	XG696 	(WX3341,WX3340);
	dff 	XG697 	(WX3343,WX3342);
	dff 	XG698 	(WX3345,WX3344);
	dff 	XG699 	(WX3347,WX3346);
	dff 	XG700 	(WX3349,WX3348);
	dff 	XG701 	(WX3351,WX3350);
	dff 	XG702 	(WX3353,WX3352);
	dff 	XG703 	(WX3355,WX3354);
	dff 	XG704 	(WX3357,WX3356);
	dff 	XG705 	(WX3359,WX3358);
	dff 	XG706 	(WX3361,WX3360);
	dff 	XG707 	(WX3363,WX3362);
	dff 	XG708 	(WX3365,WX3364);
	dff 	XG709 	(WX3367,WX3366);
	dff 	XG710 	(WX3369,WX3368);
	dff 	XG711 	(WX3371,WX3370);
	dff 	XG712 	(WX3373,WX3372);
	dff 	XG713 	(WX3375,WX3374);
	dff 	XG714 	(WX3377,WX3376);
	dff 	XG715 	(WX3379,WX3378);
	dff 	XG716 	(WX3381,WX3380);
	dff 	XG717 	(WX3383,WX3382);
	dff 	XG718 	(WX3385,WX3384);
	dff 	XG719 	(WX3387,WX3386);
	dff 	XG720 	(WX3389,WX3388);
	dff 	XG721 	(WX3391,WX3390);
	dff 	XG722 	(WX3393,WX3392);
	dff 	XG723 	(WX3395,WX3394);
	dff 	XG724 	(WX3397,WX3396);
	dff 	XG725 	(WX3399,WX3398);
	dff 	XG726 	(WX3401,WX3400);
	dff 	XG727 	(WX3403,WX3402);
	dff 	XG728 	(WX3405,WX3404);
	dff 	XG729 	(WX3407,WX3406);
	dff 	XG730 	(WX3409,WX3408);
	dff 	XG731 	(WX3411,WX3410);
	dff 	XG732 	(WX3413,WX3412);
	dff 	XG733 	(WX3415,WX3414);
	dff 	XG734 	(WX3417,WX3416);
	dff 	XG735 	(WX3419,WX3418);
	dff 	XG736 	(WX3421,WX3420);
	dff 	XG737 	(WX3423,WX3422);
	dff 	XG738 	(WX3425,WX3424);
	dff 	XG739 	(WX3427,WX3426);
	dff 	XG740 	(WX3429,WX3428);
	dff 	XG741 	(WX3431,WX3430);
	dff 	XG742 	(WX3433,WX3432);
	dff 	XG743 	(WX3435,WX3434);
	dff 	XG744 	(WX3437,WX3436);
	dff 	XG745 	(WX3439,WX3438);
	dff 	XG746 	(WX3441,WX3440);
	dff 	XG747 	(WX3443,WX3442);
	dff 	XG748 	(WX3445,WX3444);
	dff 	XG749 	(WX3447,WX3446);
	dff 	XG750 	(WX3449,WX3448);
	dff 	XG751 	(WX3451,WX3450);
	dff 	XG752 	(WX3453,WX3452);
	dff 	XG753 	(WX3455,WX3454);
	dff 	XG754 	(WX3457,WX3456);
	dff 	XG755 	(WX3459,WX3458);
	dff 	XG756 	(WX3461,WX3460);
	dff 	XG757 	(WX3463,WX3462);
	dff 	XG758 	(WX3465,WX3464);
	dff 	XG759 	(WX3467,WX3466);
	dff 	XG760 	(WX3469,WX3468);
	dff 	XG761 	(WX3471,WX3470);
	dff 	XG762 	(WX3473,WX3472);
	dff 	XG763 	(WX3475,WX3474);
	dff 	XG764 	(WX3477,WX3476);
	dff 	XG765 	(WX3479,WX3478);
	dff 	XG766 	(WX3481,WX3480);
	dff 	XG767 	(WX3483,WX3482);
	dff 	XG768 	(WX3485,WX3484);
	dff 	XG769 	(WX4364,WX4363);
	dff 	XG770 	(WX4366,WX4365);
	dff 	XG771 	(WX4368,WX4367);
	dff 	XG772 	(WX4370,WX4369);
	dff 	XG773 	(WX4372,WX4371);
	dff 	XG774 	(WX4374,WX4373);
	dff 	XG775 	(WX4376,WX4375);
	dff 	XG776 	(WX4378,WX4377);
	dff 	XG777 	(WX4380,WX4379);
	dff 	XG778 	(WX4382,WX4381);
	dff 	XG779 	(WX4384,WX4383);
	dff 	XG780 	(WX4386,WX4385);
	dff 	XG781 	(WX4388,WX4387);
	dff 	XG782 	(WX4390,WX4389);
	dff 	XG783 	(WX4392,WX4391);
	dff 	XG784 	(WX4394,WX4393);
	dff 	XG785 	(WX4396,WX4395);
	dff 	XG786 	(WX4398,WX4397);
	dff 	XG787 	(WX4400,WX4399);
	dff 	XG788 	(WX4402,WX4401);
	dff 	XG789 	(WX4404,WX4403);
	dff 	XG790 	(WX4406,WX4405);
	dff 	XG791 	(WX4408,WX4407);
	dff 	XG792 	(WX4410,WX4409);
	dff 	XG793 	(WX4412,WX4411);
	dff 	XG794 	(WX4414,WX4413);
	dff 	XG795 	(WX4416,WX4415);
	dff 	XG796 	(WX4418,WX4417);
	dff 	XG797 	(WX4420,WX4419);
	dff 	XG798 	(WX4422,WX4421);
	dff 	XG799 	(WX4424,WX4423);
	dff 	XG800 	(WX4426,WX4425);
	dff 	XG801 	(WX4524,WX4523);
	dff 	XG802 	(WX4526,WX4525);
	dff 	XG803 	(WX4528,WX4527);
	dff 	XG804 	(WX4530,WX4529);
	dff 	XG805 	(WX4532,WX4531);
	dff 	XG806 	(WX4534,WX4533);
	dff 	XG807 	(WX4536,WX4535);
	dff 	XG808 	(WX4538,WX4537);
	dff 	XG809 	(WX4540,WX4539);
	dff 	XG810 	(WX4542,WX4541);
	dff 	XG811 	(WX4544,WX4543);
	dff 	XG812 	(WX4546,WX4545);
	dff 	XG813 	(WX4548,WX4547);
	dff 	XG814 	(WX4550,WX4549);
	dff 	XG815 	(WX4552,WX4551);
	dff 	XG816 	(WX4554,WX4553);
	dff 	XG817 	(WX4556,WX4555);
	dff 	XG818 	(WX4558,WX4557);
	dff 	XG819 	(WX4560,WX4559);
	dff 	XG820 	(WX4562,WX4561);
	dff 	XG821 	(WX4564,WX4563);
	dff 	XG822 	(WX4566,WX4565);
	dff 	XG823 	(WX4568,WX4567);
	dff 	XG824 	(WX4570,WX4569);
	dff 	XG825 	(WX4572,WX4571);
	dff 	XG826 	(WX4574,WX4573);
	dff 	XG827 	(WX4576,WX4575);
	dff 	XG828 	(WX4578,WX4577);
	dff 	XG829 	(WX4580,WX4579);
	dff 	XG830 	(WX4582,WX4581);
	dff 	XG831 	(WX4584,WX4583);
	dff 	XG832 	(WX4586,WX4585);
	dff 	XG833 	(WX4588,WX4587);
	dff 	XG834 	(WX4590,WX4589);
	dff 	XG835 	(WX4592,WX4591);
	dff 	XG836 	(WX4594,WX4593);
	dff 	XG837 	(WX4596,WX4595);
	dff 	XG838 	(WX4598,WX4597);
	dff 	XG839 	(WX4600,WX4599);
	dff 	XG840 	(WX4602,WX4601);
	dff 	XG841 	(WX4604,WX4603);
	dff 	XG842 	(WX4606,WX4605);
	dff 	XG843 	(WX4608,WX4607);
	dff 	XG844 	(WX4610,WX4609);
	dff 	XG845 	(WX4612,WX4611);
	dff 	XG846 	(WX4614,WX4613);
	dff 	XG847 	(WX4616,WX4615);
	dff 	XG848 	(WX4618,WX4617);
	dff 	XG849 	(WX4620,WX4619);
	dff 	XG850 	(WX4622,WX4621);
	dff 	XG851 	(WX4624,WX4623);
	dff 	XG852 	(WX4626,WX4625);
	dff 	XG853 	(WX4628,WX4627);
	dff 	XG854 	(WX4630,WX4629);
	dff 	XG855 	(WX4632,WX4631);
	dff 	XG856 	(WX4634,WX4633);
	dff 	XG857 	(WX4636,WX4635);
	dff 	XG858 	(WX4638,WX4637);
	dff 	XG859 	(WX4640,WX4639);
	dff 	XG860 	(WX4642,WX4641);
	dff 	XG861 	(WX4644,WX4643);
	dff 	XG862 	(WX4646,WX4645);
	dff 	XG863 	(WX4648,WX4647);
	dff 	XG864 	(WX4650,WX4649);
	dff 	XG865 	(WX4652,WX4651);
	dff 	XG866 	(WX4654,WX4653);
	dff 	XG867 	(WX4656,WX4655);
	dff 	XG868 	(WX4658,WX4657);
	dff 	XG869 	(WX4660,WX4659);
	dff 	XG870 	(WX4662,WX4661);
	dff 	XG871 	(WX4664,WX4663);
	dff 	XG872 	(WX4666,WX4665);
	dff 	XG873 	(WX4668,WX4667);
	dff 	XG874 	(WX4670,WX4669);
	dff 	XG875 	(WX4672,WX4671);
	dff 	XG876 	(WX4674,WX4673);
	dff 	XG877 	(WX4676,WX4675);
	dff 	XG878 	(WX4678,WX4677);
	dff 	XG879 	(WX4680,WX4679);
	dff 	XG880 	(WX4682,WX4681);
	dff 	XG881 	(WX4684,WX4683);
	dff 	XG882 	(WX4686,WX4685);
	dff 	XG883 	(WX4688,WX4687);
	dff 	XG884 	(WX4690,WX4689);
	dff 	XG885 	(WX4692,WX4691);
	dff 	XG886 	(WX4694,WX4693);
	dff 	XG887 	(WX4696,WX4695);
	dff 	XG888 	(WX4698,WX4697);
	dff 	XG889 	(WX4700,WX4699);
	dff 	XG890 	(WX4702,WX4701);
	dff 	XG891 	(WX4704,WX4703);
	dff 	XG892 	(WX4706,WX4705);
	dff 	XG893 	(WX4708,WX4707);
	dff 	XG894 	(WX4710,WX4709);
	dff 	XG895 	(WX4712,WX4711);
	dff 	XG896 	(WX4714,WX4713);
	dff 	XG897 	(WX4716,WX4715);
	dff 	XG898 	(WX4718,WX4717);
	dff 	XG899 	(WX4720,WX4719);
	dff 	XG900 	(WX4722,WX4721);
	dff 	XG901 	(WX4724,WX4723);
	dff 	XG902 	(WX4726,WX4725);
	dff 	XG903 	(WX4728,WX4727);
	dff 	XG904 	(WX4730,WX4729);
	dff 	XG905 	(WX4732,WX4731);
	dff 	XG906 	(WX4734,WX4733);
	dff 	XG907 	(WX4736,WX4735);
	dff 	XG908 	(WX4738,WX4737);
	dff 	XG909 	(WX4740,WX4739);
	dff 	XG910 	(WX4742,WX4741);
	dff 	XG911 	(WX4744,WX4743);
	dff 	XG912 	(WX4746,WX4745);
	dff 	XG913 	(WX4748,WX4747);
	dff 	XG914 	(WX4750,WX4749);
	dff 	XG915 	(WX4752,WX4751);
	dff 	XG916 	(WX4754,WX4753);
	dff 	XG917 	(WX4756,WX4755);
	dff 	XG918 	(WX4758,WX4757);
	dff 	XG919 	(WX4760,WX4759);
	dff 	XG920 	(WX4762,WX4761);
	dff 	XG921 	(WX4764,WX4763);
	dff 	XG922 	(WX4766,WX4765);
	dff 	XG923 	(WX4768,WX4767);
	dff 	XG924 	(WX4770,WX4769);
	dff 	XG925 	(WX4772,WX4771);
	dff 	XG926 	(WX4774,WX4773);
	dff 	XG927 	(WX4776,WX4775);
	dff 	XG928 	(WX4778,WX4777);
	dff 	XG929 	(WX5657,WX5656);
	dff 	XG930 	(WX5659,WX5658);
	dff 	XG931 	(WX5661,WX5660);
	dff 	XG932 	(WX5663,WX5662);
	dff 	XG933 	(WX5665,WX5664);
	dff 	XG934 	(WX5667,WX5666);
	dff 	XG935 	(WX5669,WX5668);
	dff 	XG936 	(WX5671,WX5670);
	dff 	XG937 	(WX5673,WX5672);
	dff 	XG938 	(WX5675,WX5674);
	dff 	XG939 	(WX5677,WX5676);
	dff 	XG940 	(WX5679,WX5678);
	dff 	XG941 	(WX5681,WX5680);
	dff 	XG942 	(WX5683,WX5682);
	dff 	XG943 	(WX5685,WX5684);
	dff 	XG944 	(WX5687,WX5686);
	dff 	XG945 	(WX5689,WX5688);
	dff 	XG946 	(WX5691,WX5690);
	dff 	XG947 	(WX5693,WX5692);
	dff 	XG948 	(WX5695,WX5694);
	dff 	XG949 	(WX5697,WX5696);
	dff 	XG950 	(WX5699,WX5698);
	dff 	XG951 	(WX5701,WX5700);
	dff 	XG952 	(WX5703,WX5702);
	dff 	XG953 	(WX5705,WX5704);
	dff 	XG954 	(WX5707,WX5706);
	dff 	XG955 	(WX5709,WX5708);
	dff 	XG956 	(WX5711,WX5710);
	dff 	XG957 	(WX5713,WX5712);
	dff 	XG958 	(WX5715,WX5714);
	dff 	XG959 	(WX5717,WX5716);
	dff 	XG960 	(WX5719,WX5718);
	dff 	XG961 	(WX5817,WX5816);
	dff 	XG962 	(WX5819,WX5818);
	dff 	XG963 	(WX5821,WX5820);
	dff 	XG964 	(WX5823,WX5822);
	dff 	XG965 	(WX5825,WX5824);
	dff 	XG966 	(WX5827,WX5826);
	dff 	XG967 	(WX5829,WX5828);
	dff 	XG968 	(WX5831,WX5830);
	dff 	XG969 	(WX5833,WX5832);
	dff 	XG970 	(WX5835,WX5834);
	dff 	XG971 	(WX5837,WX5836);
	dff 	XG972 	(WX5839,WX5838);
	dff 	XG973 	(WX5841,WX5840);
	dff 	XG974 	(WX5843,WX5842);
	dff 	XG975 	(WX5845,WX5844);
	dff 	XG976 	(WX5847,WX5846);
	dff 	XG977 	(WX5849,WX5848);
	dff 	XG978 	(WX5851,WX5850);
	dff 	XG979 	(WX5853,WX5852);
	dff 	XG980 	(WX5855,WX5854);
	dff 	XG981 	(WX5857,WX5856);
	dff 	XG982 	(WX5859,WX5858);
	dff 	XG983 	(WX5861,WX5860);
	dff 	XG984 	(WX5863,WX5862);
	dff 	XG985 	(WX5865,WX5864);
	dff 	XG986 	(WX5867,WX5866);
	dff 	XG987 	(WX5869,WX5868);
	dff 	XG988 	(WX5871,WX5870);
	dff 	XG989 	(WX5873,WX5872);
	dff 	XG990 	(WX5875,WX5874);
	dff 	XG991 	(WX5877,WX5876);
	dff 	XG992 	(WX5879,WX5878);
	dff 	XG993 	(WX5881,WX5880);
	dff 	XG994 	(WX5883,WX5882);
	dff 	XG995 	(WX5885,WX5884);
	dff 	XG996 	(WX5887,WX5886);
	dff 	XG997 	(WX5889,WX5888);
	dff 	XG998 	(WX5891,WX5890);
	dff 	XG999 	(WX5893,WX5892);
	dff 	XG1000 	(WX5895,WX5894);
	dff 	XG1001 	(WX5897,WX5896);
	dff 	XG1002 	(WX5899,WX5898);
	dff 	XG1003 	(WX5901,WX5900);
	dff 	XG1004 	(WX5903,WX5902);
	dff 	XG1005 	(WX5905,WX5904);
	dff 	XG1006 	(WX5907,WX5906);
	dff 	XG1007 	(WX5909,WX5908);
	dff 	XG1008 	(WX5911,WX5910);
	dff 	XG1009 	(WX5913,WX5912);
	dff 	XG1010 	(WX5915,WX5914);
	dff 	XG1011 	(WX5917,WX5916);
	dff 	XG1012 	(WX5919,WX5918);
	dff 	XG1013 	(WX5921,WX5920);
	dff 	XG1014 	(WX5923,WX5922);
	dff 	XG1015 	(WX5925,WX5924);
	dff 	XG1016 	(WX5927,WX5926);
	dff 	XG1017 	(WX5929,WX5928);
	dff 	XG1018 	(WX5931,WX5930);
	dff 	XG1019 	(WX5933,WX5932);
	dff 	XG1020 	(WX5935,WX5934);
	dff 	XG1021 	(WX5937,WX5936);
	dff 	XG1022 	(WX5939,WX5938);
	dff 	XG1023 	(WX5941,WX5940);
	dff 	XG1024 	(WX5943,WX5942);
	dff 	XG1025 	(WX5945,WX5944);
	dff 	XG1026 	(WX5947,WX5946);
	dff 	XG1027 	(WX5949,WX5948);
	dff 	XG1028 	(WX5951,WX5950);
	dff 	XG1029 	(WX5953,WX5952);
	dff 	XG1030 	(WX5955,WX5954);
	dff 	XG1031 	(WX5957,WX5956);
	dff 	XG1032 	(WX5959,WX5958);
	dff 	XG1033 	(WX5961,WX5960);
	dff 	XG1034 	(WX5963,WX5962);
	dff 	XG1035 	(WX5965,WX5964);
	dff 	XG1036 	(WX5967,WX5966);
	dff 	XG1037 	(WX5969,WX5968);
	dff 	XG1038 	(WX5971,WX5970);
	dff 	XG1039 	(WX5973,WX5972);
	dff 	XG1040 	(WX5975,WX5974);
	dff 	XG1041 	(WX5977,WX5976);
	dff 	XG1042 	(WX5979,WX5978);
	dff 	XG1043 	(WX5981,WX5980);
	dff 	XG1044 	(WX5983,WX5982);
	dff 	XG1045 	(WX5985,WX5984);
	dff 	XG1046 	(WX5987,WX5986);
	dff 	XG1047 	(WX5989,WX5988);
	dff 	XG1048 	(WX5991,WX5990);
	dff 	XG1049 	(WX5993,WX5992);
	dff 	XG1050 	(WX5995,WX5994);
	dff 	XG1051 	(WX5997,WX5996);
	dff 	XG1052 	(WX5999,WX5998);
	dff 	XG1053 	(WX6001,WX6000);
	dff 	XG1054 	(WX6003,WX6002);
	dff 	XG1055 	(WX6005,WX6004);
	dff 	XG1056 	(WX6007,WX6006);
	dff 	XG1057 	(WX6009,WX6008);
	dff 	XG1058 	(WX6011,WX6010);
	dff 	XG1059 	(WX6013,WX6012);
	dff 	XG1060 	(WX6015,WX6014);
	dff 	XG1061 	(WX6017,WX6016);
	dff 	XG1062 	(WX6019,WX6018);
	dff 	XG1063 	(WX6021,WX6020);
	dff 	XG1064 	(WX6023,WX6022);
	dff 	XG1065 	(WX6025,WX6024);
	dff 	XG1066 	(WX6027,WX6026);
	dff 	XG1067 	(WX6029,WX6028);
	dff 	XG1068 	(WX6031,WX6030);
	dff 	XG1069 	(WX6033,WX6032);
	dff 	XG1070 	(WX6035,WX6034);
	dff 	XG1071 	(WX6037,WX6036);
	dff 	XG1072 	(WX6039,WX6038);
	dff 	XG1073 	(WX6041,WX6040);
	dff 	XG1074 	(WX6043,WX6042);
	dff 	XG1075 	(WX6045,WX6044);
	dff 	XG1076 	(WX6047,WX6046);
	dff 	XG1077 	(WX6049,WX6048);
	dff 	XG1078 	(WX6051,WX6050);
	dff 	XG1079 	(WX6053,WX6052);
	dff 	XG1080 	(WX6055,WX6054);
	dff 	XG1081 	(WX6057,WX6056);
	dff 	XG1082 	(WX6059,WX6058);
	dff 	XG1083 	(WX6061,WX6060);
	dff 	XG1084 	(WX6063,WX6062);
	dff 	XG1085 	(WX6065,WX6064);
	dff 	XG1086 	(WX6067,WX6066);
	dff 	XG1087 	(WX6069,WX6068);
	dff 	XG1088 	(WX6071,WX6070);
	dff 	XG1089 	(WX6950,WX6949);
	dff 	XG1090 	(WX6952,WX6951);
	dff 	XG1091 	(WX6954,WX6953);
	dff 	XG1092 	(WX6956,WX6955);
	dff 	XG1093 	(WX6958,WX6957);
	dff 	XG1094 	(WX6960,WX6959);
	dff 	XG1095 	(WX6962,WX6961);
	dff 	XG1096 	(WX6964,WX6963);
	dff 	XG1097 	(WX6966,WX6965);
	dff 	XG1098 	(WX6968,WX6967);
	dff 	XG1099 	(WX6970,WX6969);
	dff 	XG1100 	(WX6972,WX6971);
	dff 	XG1101 	(WX6974,WX6973);
	dff 	XG1102 	(WX6976,WX6975);
	dff 	XG1103 	(WX6978,WX6977);
	dff 	XG1104 	(WX6980,WX6979);
	dff 	XG1105 	(WX6982,WX6981);
	dff 	XG1106 	(WX6984,WX6983);
	dff 	XG1107 	(WX6986,WX6985);
	dff 	XG1108 	(WX6988,WX6987);
	dff 	XG1109 	(WX6990,WX6989);
	dff 	XG1110 	(WX6992,WX6991);
	dff 	XG1111 	(WX6994,WX6993);
	dff 	XG1112 	(WX6996,WX6995);
	dff 	XG1113 	(WX6998,WX6997);
	dff 	XG1114 	(WX7000,WX6999);
	dff 	XG1115 	(WX7002,WX7001);
	dff 	XG1116 	(WX7004,WX7003);
	dff 	XG1117 	(WX7006,WX7005);
	dff 	XG1118 	(WX7008,WX7007);
	dff 	XG1119 	(WX7010,WX7009);
	dff 	XG1120 	(WX7012,WX7011);
	dff 	XG1121 	(WX7110,WX7109);
	dff 	XG1122 	(WX7112,WX7111);
	dff 	XG1123 	(WX7114,WX7113);
	dff 	XG1124 	(WX7116,WX7115);
	dff 	XG1125 	(WX7118,WX7117);
	dff 	XG1126 	(WX7120,WX7119);
	dff 	XG1127 	(WX7122,WX7121);
	dff 	XG1128 	(WX7124,WX7123);
	dff 	XG1129 	(WX7126,WX7125);
	dff 	XG1130 	(WX7128,WX7127);
	dff 	XG1131 	(WX7130,WX7129);
	dff 	XG1132 	(WX7132,WX7131);
	dff 	XG1133 	(WX7134,WX7133);
	dff 	XG1134 	(WX7136,WX7135);
	dff 	XG1135 	(WX7138,WX7137);
	dff 	XG1136 	(WX7140,WX7139);
	dff 	XG1137 	(WX7142,WX7141);
	dff 	XG1138 	(WX7144,WX7143);
	dff 	XG1139 	(WX7146,WX7145);
	dff 	XG1140 	(WX7148,WX7147);
	dff 	XG1141 	(WX7150,WX7149);
	dff 	XG1142 	(WX7152,WX7151);
	dff 	XG1143 	(WX7154,WX7153);
	dff 	XG1144 	(WX7156,WX7155);
	dff 	XG1145 	(WX7158,WX7157);
	dff 	XG1146 	(WX7160,WX7159);
	dff 	XG1147 	(WX7162,WX7161);
	dff 	XG1148 	(WX7164,WX7163);
	dff 	XG1149 	(WX7166,WX7165);
	dff 	XG1150 	(WX7168,WX7167);
	dff 	XG1151 	(WX7170,WX7169);
	dff 	XG1152 	(WX7172,WX7171);
	dff 	XG1153 	(WX7174,WX7173);
	dff 	XG1154 	(WX7176,WX7175);
	dff 	XG1155 	(WX7178,WX7177);
	dff 	XG1156 	(WX7180,WX7179);
	dff 	XG1157 	(WX7182,WX7181);
	dff 	XG1158 	(WX7184,WX7183);
	dff 	XG1159 	(WX7186,WX7185);
	dff 	XG1160 	(WX7188,WX7187);
	dff 	XG1161 	(WX7190,WX7189);
	dff 	XG1162 	(WX7192,WX7191);
	dff 	XG1163 	(WX7194,WX7193);
	dff 	XG1164 	(WX7196,WX7195);
	dff 	XG1165 	(WX7198,WX7197);
	dff 	XG1166 	(WX7200,WX7199);
	dff 	XG1167 	(WX7202,WX7201);
	dff 	XG1168 	(WX7204,WX7203);
	dff 	XG1169 	(WX7206,WX7205);
	dff 	XG1170 	(WX7208,WX7207);
	dff 	XG1171 	(WX7210,WX7209);
	dff 	XG1172 	(WX7212,WX7211);
	dff 	XG1173 	(WX7214,WX7213);
	dff 	XG1174 	(WX7216,WX7215);
	dff 	XG1175 	(WX7218,WX7217);
	dff 	XG1176 	(WX7220,WX7219);
	dff 	XG1177 	(WX7222,WX7221);
	dff 	XG1178 	(WX7224,WX7223);
	dff 	XG1179 	(WX7226,WX7225);
	dff 	XG1180 	(WX7228,WX7227);
	dff 	XG1181 	(WX7230,WX7229);
	dff 	XG1182 	(WX7232,WX7231);
	dff 	XG1183 	(WX7234,WX7233);
	dff 	XG1184 	(WX7236,WX7235);
	dff 	XG1185 	(WX7238,WX7237);
	dff 	XG1186 	(WX7240,WX7239);
	dff 	XG1187 	(WX7242,WX7241);
	dff 	XG1188 	(WX7244,WX7243);
	dff 	XG1189 	(WX7246,WX7245);
	dff 	XG1190 	(WX7248,WX7247);
	dff 	XG1191 	(WX7250,WX7249);
	dff 	XG1192 	(WX7252,WX7251);
	dff 	XG1193 	(WX7254,WX7253);
	dff 	XG1194 	(WX7256,WX7255);
	dff 	XG1195 	(WX7258,WX7257);
	dff 	XG1196 	(WX7260,WX7259);
	dff 	XG1197 	(WX7262,WX7261);
	dff 	XG1198 	(WX7264,WX7263);
	dff 	XG1199 	(WX7266,WX7265);
	dff 	XG1200 	(WX7268,WX7267);
	dff 	XG1201 	(WX7270,WX7269);
	dff 	XG1202 	(WX7272,WX7271);
	dff 	XG1203 	(WX7274,WX7273);
	dff 	XG1204 	(WX7276,WX7275);
	dff 	XG1205 	(WX7278,WX7277);
	dff 	XG1206 	(WX7280,WX7279);
	dff 	XG1207 	(WX7282,WX7281);
	dff 	XG1208 	(WX7284,WX7283);
	dff 	XG1209 	(WX7286,WX7285);
	dff 	XG1210 	(WX7288,WX7287);
	dff 	XG1211 	(WX7290,WX7289);
	dff 	XG1212 	(WX7292,WX7291);
	dff 	XG1213 	(WX7294,WX7293);
	dff 	XG1214 	(WX7296,WX7295);
	dff 	XG1215 	(WX7298,WX7297);
	dff 	XG1216 	(WX7300,WX7299);
	dff 	XG1217 	(WX7302,WX7301);
	dff 	XG1218 	(WX7304,WX7303);
	dff 	XG1219 	(WX7306,WX7305);
	dff 	XG1220 	(WX7308,WX7307);
	dff 	XG1221 	(WX7310,WX7309);
	dff 	XG1222 	(WX7312,WX7311);
	dff 	XG1223 	(WX7314,WX7313);
	dff 	XG1224 	(WX7316,WX7315);
	dff 	XG1225 	(WX7318,WX7317);
	dff 	XG1226 	(WX7320,WX7319);
	dff 	XG1227 	(WX7322,WX7321);
	dff 	XG1228 	(WX7324,WX7323);
	dff 	XG1229 	(WX7326,WX7325);
	dff 	XG1230 	(WX7328,WX7327);
	dff 	XG1231 	(WX7330,WX7329);
	dff 	XG1232 	(WX7332,WX7331);
	dff 	XG1233 	(WX7334,WX7333);
	dff 	XG1234 	(WX7336,WX7335);
	dff 	XG1235 	(WX7338,WX7337);
	dff 	XG1236 	(WX7340,WX7339);
	dff 	XG1237 	(WX7342,WX7341);
	dff 	XG1238 	(WX7344,WX7343);
	dff 	XG1239 	(WX7346,WX7345);
	dff 	XG1240 	(WX7348,WX7347);
	dff 	XG1241 	(WX7350,WX7349);
	dff 	XG1242 	(WX7352,WX7351);
	dff 	XG1243 	(WX7354,WX7353);
	dff 	XG1244 	(WX7356,WX7355);
	dff 	XG1245 	(WX7358,WX7357);
	dff 	XG1246 	(WX7360,WX7359);
	dff 	XG1247 	(WX7362,WX7361);
	dff 	XG1248 	(WX7364,WX7363);
	dff 	XG1249 	(WX8243,WX8242);
	dff 	XG1250 	(WX8245,WX8244);
	dff 	XG1251 	(WX8247,WX8246);
	dff 	XG1252 	(WX8249,WX8248);
	dff 	XG1253 	(WX8251,WX8250);
	dff 	XG1254 	(WX8253,WX8252);
	dff 	XG1255 	(WX8255,WX8254);
	dff 	XG1256 	(WX8257,WX8256);
	dff 	XG1257 	(WX8259,WX8258);
	dff 	XG1258 	(WX8261,WX8260);
	dff 	XG1259 	(WX8263,WX8262);
	dff 	XG1260 	(WX8265,WX8264);
	dff 	XG1261 	(WX8267,WX8266);
	dff 	XG1262 	(WX8269,WX8268);
	dff 	XG1263 	(WX8271,WX8270);
	dff 	XG1264 	(WX8273,WX8272);
	dff 	XG1265 	(WX8275,WX8274);
	dff 	XG1266 	(WX8277,WX8276);
	dff 	XG1267 	(WX8279,WX8278);
	dff 	XG1268 	(WX8281,WX8280);
	dff 	XG1269 	(WX8283,WX8282);
	dff 	XG1270 	(WX8285,WX8284);
	dff 	XG1271 	(WX8287,WX8286);
	dff 	XG1272 	(WX8289,WX8288);
	dff 	XG1273 	(WX8291,WX8290);
	dff 	XG1274 	(WX8293,WX8292);
	dff 	XG1275 	(WX8295,WX8294);
	dff 	XG1276 	(WX8297,WX8296);
	dff 	XG1277 	(WX8299,WX8298);
	dff 	XG1278 	(WX8301,WX8300);
	dff 	XG1279 	(WX8303,WX8302);
	dff 	XG1280 	(WX8305,WX8304);
	dff 	XG1281 	(WX8403,WX8402);
	dff 	XG1282 	(WX8405,WX8404);
	dff 	XG1283 	(WX8407,WX8406);
	dff 	XG1284 	(WX8409,WX8408);
	dff 	XG1285 	(WX8411,WX8410);
	dff 	XG1286 	(WX8413,WX8412);
	dff 	XG1287 	(WX8415,WX8414);
	dff 	XG1288 	(WX8417,WX8416);
	dff 	XG1289 	(WX8419,WX8418);
	dff 	XG1290 	(WX8421,WX8420);
	dff 	XG1291 	(WX8423,WX8422);
	dff 	XG1292 	(WX8425,WX8424);
	dff 	XG1293 	(WX8427,WX8426);
	dff 	XG1294 	(WX8429,WX8428);
	dff 	XG1295 	(WX8431,WX8430);
	dff 	XG1296 	(WX8433,WX8432);
	dff 	XG1297 	(WX8435,WX8434);
	dff 	XG1298 	(WX8437,WX8436);
	dff 	XG1299 	(WX8439,WX8438);
	dff 	XG1300 	(WX8441,WX8440);
	dff 	XG1301 	(WX8443,WX8442);
	dff 	XG1302 	(WX8445,WX8444);
	dff 	XG1303 	(WX8447,WX8446);
	dff 	XG1304 	(WX8449,WX8448);
	dff 	XG1305 	(WX8451,WX8450);
	dff 	XG1306 	(WX8453,WX8452);
	dff 	XG1307 	(WX8455,WX8454);
	dff 	XG1308 	(WX8457,WX8456);
	dff 	XG1309 	(WX8459,WX8458);
	dff 	XG1310 	(WX8461,WX8460);
	dff 	XG1311 	(WX8463,WX8462);
	dff 	XG1312 	(WX8465,WX8464);
	dff 	XG1313 	(WX8467,WX8466);
	dff 	XG1314 	(WX8469,WX8468);
	dff 	XG1315 	(WX8471,WX8470);
	dff 	XG1316 	(WX8473,WX8472);
	dff 	XG1317 	(WX8475,WX8474);
	dff 	XG1318 	(WX8477,WX8476);
	dff 	XG1319 	(WX8479,WX8478);
	dff 	XG1320 	(WX8481,WX8480);
	dff 	XG1321 	(WX8483,WX8482);
	dff 	XG1322 	(WX8485,WX8484);
	dff 	XG1323 	(WX8487,WX8486);
	dff 	XG1324 	(WX8489,WX8488);
	dff 	XG1325 	(WX8491,WX8490);
	dff 	XG1326 	(WX8493,WX8492);
	dff 	XG1327 	(WX8495,WX8494);
	dff 	XG1328 	(WX8497,WX8496);
	dff 	XG1329 	(WX8499,WX8498);
	dff 	XG1330 	(WX8501,WX8500);
	dff 	XG1331 	(WX8503,WX8502);
	dff 	XG1332 	(WX8505,WX8504);
	dff 	XG1333 	(WX8507,WX8506);
	dff 	XG1334 	(WX8509,WX8508);
	dff 	XG1335 	(WX8511,WX8510);
	dff 	XG1336 	(WX8513,WX8512);
	dff 	XG1337 	(WX8515,WX8514);
	dff 	XG1338 	(WX8517,WX8516);
	dff 	XG1339 	(WX8519,WX8518);
	dff 	XG1340 	(WX8521,WX8520);
	dff 	XG1341 	(WX8523,WX8522);
	dff 	XG1342 	(WX8525,WX8524);
	dff 	XG1343 	(WX8527,WX8526);
	dff 	XG1344 	(WX8529,WX8528);
	dff 	XG1345 	(WX8531,WX8530);
	dff 	XG1346 	(WX8533,WX8532);
	dff 	XG1347 	(WX8535,WX8534);
	dff 	XG1348 	(WX8537,WX8536);
	dff 	XG1349 	(WX8539,WX8538);
	dff 	XG1350 	(WX8541,WX8540);
	dff 	XG1351 	(WX8543,WX8542);
	dff 	XG1352 	(WX8545,WX8544);
	dff 	XG1353 	(WX8547,WX8546);
	dff 	XG1354 	(WX8549,WX8548);
	dff 	XG1355 	(WX8551,WX8550);
	dff 	XG1356 	(WX8553,WX8552);
	dff 	XG1357 	(WX8555,WX8554);
	dff 	XG1358 	(WX8557,WX8556);
	dff 	XG1359 	(WX8559,WX8558);
	dff 	XG1360 	(WX8561,WX8560);
	dff 	XG1361 	(WX8563,WX8562);
	dff 	XG1362 	(WX8565,WX8564);
	dff 	XG1363 	(WX8567,WX8566);
	dff 	XG1364 	(WX8569,WX8568);
	dff 	XG1365 	(WX8571,WX8570);
	dff 	XG1366 	(WX8573,WX8572);
	dff 	XG1367 	(WX8575,WX8574);
	dff 	XG1368 	(WX8577,WX8576);
	dff 	XG1369 	(WX8579,WX8578);
	dff 	XG1370 	(WX8581,WX8580);
	dff 	XG1371 	(WX8583,WX8582);
	dff 	XG1372 	(WX8585,WX8584);
	dff 	XG1373 	(WX8587,WX8586);
	dff 	XG1374 	(WX8589,WX8588);
	dff 	XG1375 	(WX8591,WX8590);
	dff 	XG1376 	(WX8593,WX8592);
	dff 	XG1377 	(WX8595,WX8594);
	dff 	XG1378 	(WX8597,WX8596);
	dff 	XG1379 	(WX8599,WX8598);
	dff 	XG1380 	(WX8601,WX8600);
	dff 	XG1381 	(WX8603,WX8602);
	dff 	XG1382 	(WX8605,WX8604);
	dff 	XG1383 	(WX8607,WX8606);
	dff 	XG1384 	(WX8609,WX8608);
	dff 	XG1385 	(WX8611,WX8610);
	dff 	XG1386 	(WX8613,WX8612);
	dff 	XG1387 	(WX8615,WX8614);
	dff 	XG1388 	(WX8617,WX8616);
	dff 	XG1389 	(WX8619,WX8618);
	dff 	XG1390 	(WX8621,WX8620);
	dff 	XG1391 	(WX8623,WX8622);
	dff 	XG1392 	(WX8625,WX8624);
	dff 	XG1393 	(WX8627,WX8626);
	dff 	XG1394 	(WX8629,WX8628);
	dff 	XG1395 	(WX8631,WX8630);
	dff 	XG1396 	(WX8633,WX8632);
	dff 	XG1397 	(WX8635,WX8634);
	dff 	XG1398 	(WX8637,WX8636);
	dff 	XG1399 	(WX8639,WX8638);
	dff 	XG1400 	(WX8641,WX8640);
	dff 	XG1401 	(WX8643,WX8642);
	dff 	XG1402 	(WX8645,WX8644);
	dff 	XG1403 	(WX8647,WX8646);
	dff 	XG1404 	(WX8649,WX8648);
	dff 	XG1405 	(WX8651,WX8650);
	dff 	XG1406 	(WX8653,WX8652);
	dff 	XG1407 	(WX8655,WX8654);
	dff 	XG1408 	(WX8657,WX8656);
	dff 	XG1409 	(WX9536,WX9535);
	dff 	XG1410 	(WX9538,WX9537);
	dff 	XG1411 	(WX9540,WX9539);
	dff 	XG1412 	(WX9542,WX9541);
	dff 	XG1413 	(WX9544,WX9543);
	dff 	XG1414 	(WX9546,WX9545);
	dff 	XG1415 	(WX9548,WX9547);
	dff 	XG1416 	(WX9550,WX9549);
	dff 	XG1417 	(WX9552,WX9551);
	dff 	XG1418 	(WX9554,WX9553);
	dff 	XG1419 	(WX9556,WX9555);
	dff 	XG1420 	(WX9558,WX9557);
	dff 	XG1421 	(WX9560,WX9559);
	dff 	XG1422 	(WX9562,WX9561);
	dff 	XG1423 	(WX9564,WX9563);
	dff 	XG1424 	(WX9566,WX9565);
	dff 	XG1425 	(WX9568,WX9567);
	dff 	XG1426 	(WX9570,WX9569);
	dff 	XG1427 	(WX9572,WX9571);
	dff 	XG1428 	(WX9574,WX9573);
	dff 	XG1429 	(WX9576,WX9575);
	dff 	XG1430 	(WX9578,WX9577);
	dff 	XG1431 	(WX9580,WX9579);
	dff 	XG1432 	(WX9582,WX9581);
	dff 	XG1433 	(WX9584,WX9583);
	dff 	XG1434 	(WX9586,WX9585);
	dff 	XG1435 	(WX9588,WX9587);
	dff 	XG1436 	(WX9590,WX9589);
	dff 	XG1437 	(WX9592,WX9591);
	dff 	XG1438 	(WX9594,WX9593);
	dff 	XG1439 	(WX9596,WX9595);
	dff 	XG1440 	(WX9598,WX9597);
	dff 	XG1441 	(WX9696,WX9695);
	dff 	XG1442 	(WX9698,WX9697);
	dff 	XG1443 	(WX9700,WX9699);
	dff 	XG1444 	(WX9702,WX9701);
	dff 	XG1445 	(WX9704,WX9703);
	dff 	XG1446 	(WX9706,WX9705);
	dff 	XG1447 	(WX9708,WX9707);
	dff 	XG1448 	(WX9710,WX9709);
	dff 	XG1449 	(WX9712,WX9711);
	dff 	XG1450 	(WX9714,WX9713);
	dff 	XG1451 	(WX9716,WX9715);
	dff 	XG1452 	(WX9718,WX9717);
	dff 	XG1453 	(WX9720,WX9719);
	dff 	XG1454 	(WX9722,WX9721);
	dff 	XG1455 	(WX9724,WX9723);
	dff 	XG1456 	(WX9726,WX9725);
	dff 	XG1457 	(WX9728,WX9727);
	dff 	XG1458 	(WX9730,WX9729);
	dff 	XG1459 	(WX9732,WX9731);
	dff 	XG1460 	(WX9734,WX9733);
	dff 	XG1461 	(WX9736,WX9735);
	dff 	XG1462 	(WX9738,WX9737);
	dff 	XG1463 	(WX9740,WX9739);
	dff 	XG1464 	(WX9742,WX9741);
	dff 	XG1465 	(WX9744,WX9743);
	dff 	XG1466 	(WX9746,WX9745);
	dff 	XG1467 	(WX9748,WX9747);
	dff 	XG1468 	(WX9750,WX9749);
	dff 	XG1469 	(WX9752,WX9751);
	dff 	XG1470 	(WX9754,WX9753);
	dff 	XG1471 	(WX9756,WX9755);
	dff 	XG1472 	(WX9758,WX9757);
	dff 	XG1473 	(WX9760,WX9759);
	dff 	XG1474 	(WX9762,WX9761);
	dff 	XG1475 	(WX9764,WX9763);
	dff 	XG1476 	(WX9766,WX9765);
	dff 	XG1477 	(WX9768,WX9767);
	dff 	XG1478 	(WX9770,WX9769);
	dff 	XG1479 	(WX9772,WX9771);
	dff 	XG1480 	(WX9774,WX9773);
	dff 	XG1481 	(WX9776,WX9775);
	dff 	XG1482 	(WX9778,WX9777);
	dff 	XG1483 	(WX9780,WX9779);
	dff 	XG1484 	(WX9782,WX9781);
	dff 	XG1485 	(WX9784,WX9783);
	dff 	XG1486 	(WX9786,WX9785);
	dff 	XG1487 	(WX9788,WX9787);
	dff 	XG1488 	(WX9790,WX9789);
	dff 	XG1489 	(WX9792,WX9791);
	dff 	XG1490 	(WX9794,WX9793);
	dff 	XG1491 	(WX9796,WX9795);
	dff 	XG1492 	(WX9798,WX9797);
	dff 	XG1493 	(WX9800,WX9799);
	dff 	XG1494 	(WX9802,WX9801);
	dff 	XG1495 	(WX9804,WX9803);
	dff 	XG1496 	(WX9806,WX9805);
	dff 	XG1497 	(WX9808,WX9807);
	dff 	XG1498 	(WX9810,WX9809);
	dff 	XG1499 	(WX9812,WX9811);
	dff 	XG1500 	(WX9814,WX9813);
	dff 	XG1501 	(WX9816,WX9815);
	dff 	XG1502 	(WX9818,WX9817);
	dff 	XG1503 	(WX9820,WX9819);
	dff 	XG1504 	(WX9822,WX9821);
	dff 	XG1505 	(WX9824,WX9823);
	dff 	XG1506 	(WX9826,WX9825);
	dff 	XG1507 	(WX9828,WX9827);
	dff 	XG1508 	(WX9830,WX9829);
	dff 	XG1509 	(WX9832,WX9831);
	dff 	XG1510 	(WX9834,WX9833);
	dff 	XG1511 	(WX9836,WX9835);
	dff 	XG1512 	(WX9838,WX9837);
	dff 	XG1513 	(WX9840,WX9839);
	dff 	XG1514 	(WX9842,WX9841);
	dff 	XG1515 	(WX9844,WX9843);
	dff 	XG1516 	(WX9846,WX9845);
	dff 	XG1517 	(WX9848,WX9847);
	dff 	XG1518 	(WX9850,WX9849);
	dff 	XG1519 	(WX9852,WX9851);
	dff 	XG1520 	(WX9854,WX9853);
	dff 	XG1521 	(WX9856,WX9855);
	dff 	XG1522 	(WX9858,WX9857);
	dff 	XG1523 	(WX9860,WX9859);
	dff 	XG1524 	(WX9862,WX9861);
	dff 	XG1525 	(WX9864,WX9863);
	dff 	XG1526 	(WX9866,WX9865);
	dff 	XG1527 	(WX9868,WX9867);
	dff 	XG1528 	(WX9870,WX9869);
	dff 	XG1529 	(WX9872,WX9871);
	dff 	XG1530 	(WX9874,WX9873);
	dff 	XG1531 	(WX9876,WX9875);
	dff 	XG1532 	(WX9878,WX9877);
	dff 	XG1533 	(WX9880,WX9879);
	dff 	XG1534 	(WX9882,WX9881);
	dff 	XG1535 	(WX9884,WX9883);
	dff 	XG1536 	(WX9886,WX9885);
	dff 	XG1537 	(WX9888,WX9887);
	dff 	XG1538 	(WX9890,WX9889);
	dff 	XG1539 	(WX9892,WX9891);
	dff 	XG1540 	(WX9894,WX9893);
	dff 	XG1541 	(WX9896,WX9895);
	dff 	XG1542 	(WX9898,WX9897);
	dff 	XG1543 	(WX9900,WX9899);
	dff 	XG1544 	(WX9902,WX9901);
	dff 	XG1545 	(WX9904,WX9903);
	dff 	XG1546 	(WX9906,WX9905);
	dff 	XG1547 	(WX9908,WX9907);
	dff 	XG1548 	(WX9910,WX9909);
	dff 	XG1549 	(WX9912,WX9911);
	dff 	XG1550 	(WX9914,WX9913);
	dff 	XG1551 	(WX9916,WX9915);
	dff 	XG1552 	(WX9918,WX9917);
	dff 	XG1553 	(WX9920,WX9919);
	dff 	XG1554 	(WX9922,WX9921);
	dff 	XG1555 	(WX9924,WX9923);
	dff 	XG1556 	(WX9926,WX9925);
	dff 	XG1557 	(WX9928,WX9927);
	dff 	XG1558 	(WX9930,WX9929);
	dff 	XG1559 	(WX9932,WX9931);
	dff 	XG1560 	(WX9934,WX9933);
	dff 	XG1561 	(WX9936,WX9935);
	dff 	XG1562 	(WX9938,WX9937);
	dff 	XG1563 	(WX9940,WX9939);
	dff 	XG1564 	(WX9942,WX9941);
	dff 	XG1565 	(WX9944,WX9943);
	dff 	XG1566 	(WX9946,WX9945);
	dff 	XG1567 	(WX9948,WX9947);
	dff 	XG1568 	(WX9950,WX9949);
	dff 	XG1569 	(WX10829,WX10828);
	dff 	XG1570 	(WX10831,WX10830);
	dff 	XG1571 	(WX10833,WX10832);
	dff 	XG1572 	(WX10835,WX10834);
	dff 	XG1573 	(WX10837,WX10836);
	dff 	XG1574 	(WX10839,WX10838);
	dff 	XG1575 	(WX10841,WX10840);
	dff 	XG1576 	(WX10843,WX10842);
	dff 	XG1577 	(WX10845,WX10844);
	dff 	XG1578 	(WX10847,WX10846);
	dff 	XG1579 	(WX10849,WX10848);
	dff 	XG1580 	(WX10851,WX10850);
	dff 	XG1581 	(WX10853,WX10852);
	dff 	XG1582 	(WX10855,WX10854);
	dff 	XG1583 	(WX10857,WX10856);
	dff 	XG1584 	(WX10859,WX10858);
	dff 	XG1585 	(WX10861,WX10860);
	dff 	XG1586 	(WX10863,WX10862);
	dff 	XG1587 	(WX10865,WX10864);
	dff 	XG1588 	(WX10867,WX10866);
	dff 	XG1589 	(WX10869,WX10868);
	dff 	XG1590 	(WX10871,WX10870);
	dff 	XG1591 	(WX10873,WX10872);
	dff 	XG1592 	(WX10875,WX10874);
	dff 	XG1593 	(WX10877,WX10876);
	dff 	XG1594 	(WX10879,WX10878);
	dff 	XG1595 	(WX10881,WX10880);
	dff 	XG1596 	(WX10883,WX10882);
	dff 	XG1597 	(WX10885,WX10884);
	dff 	XG1598 	(WX10887,WX10886);
	dff 	XG1599 	(WX10889,WX10888);
	dff 	XG1600 	(WX10891,WX10890);
	dff 	XG1601 	(WX10989,WX10988);
	dff 	XG1602 	(WX10991,WX10990);
	dff 	XG1603 	(WX10993,WX10992);
	dff 	XG1604 	(WX10995,WX10994);
	dff 	XG1605 	(WX10997,WX10996);
	dff 	XG1606 	(WX10999,WX10998);
	dff 	XG1607 	(WX11001,WX11000);
	dff 	XG1608 	(WX11003,WX11002);
	dff 	XG1609 	(WX11005,WX11004);
	dff 	XG1610 	(WX11007,WX11006);
	dff 	XG1611 	(WX11009,WX11008);
	dff 	XG1612 	(WX11011,WX11010);
	dff 	XG1613 	(WX11013,WX11012);
	dff 	XG1614 	(WX11015,WX11014);
	dff 	XG1615 	(WX11017,WX11016);
	dff 	XG1616 	(WX11019,WX11018);
	dff 	XG1617 	(WX11021,WX11020);
	dff 	XG1618 	(WX11023,WX11022);
	dff 	XG1619 	(WX11025,WX11024);
	dff 	XG1620 	(WX11027,WX11026);
	dff 	XG1621 	(WX11029,WX11028);
	dff 	XG1622 	(WX11031,WX11030);
	dff 	XG1623 	(WX11033,WX11032);
	dff 	XG1624 	(WX11035,WX11034);
	dff 	XG1625 	(WX11037,WX11036);
	dff 	XG1626 	(WX11039,WX11038);
	dff 	XG1627 	(WX11041,WX11040);
	dff 	XG1628 	(WX11043,WX11042);
	dff 	XG1629 	(WX11045,WX11044);
	dff 	XG1630 	(WX11047,WX11046);
	dff 	XG1631 	(WX11049,WX11048);
	dff 	XG1632 	(WX11051,WX11050);
	dff 	XG1633 	(WX11053,WX11052);
	dff 	XG1634 	(WX11055,WX11054);
	dff 	XG1635 	(WX11057,WX11056);
	dff 	XG1636 	(WX11059,WX11058);
	dff 	XG1637 	(WX11061,WX11060);
	dff 	XG1638 	(WX11063,WX11062);
	dff 	XG1639 	(WX11065,WX11064);
	dff 	XG1640 	(WX11067,WX11066);
	dff 	XG1641 	(WX11069,WX11068);
	dff 	XG1642 	(WX11071,WX11070);
	dff 	XG1643 	(WX11073,WX11072);
	dff 	XG1644 	(WX11075,WX11074);
	dff 	XG1645 	(WX11077,WX11076);
	dff 	XG1646 	(WX11079,WX11078);
	dff 	XG1647 	(WX11081,WX11080);
	dff 	XG1648 	(WX11083,WX11082);
	dff 	XG1649 	(WX11085,WX11084);
	dff 	XG1650 	(WX11087,WX11086);
	dff 	XG1651 	(WX11089,WX11088);
	dff 	XG1652 	(WX11091,WX11090);
	dff 	XG1653 	(WX11093,WX11092);
	dff 	XG1654 	(WX11095,WX11094);
	dff 	XG1655 	(WX11097,WX11096);
	dff 	XG1656 	(WX11099,WX11098);
	dff 	XG1657 	(WX11101,WX11100);
	dff 	XG1658 	(WX11103,WX11102);
	dff 	XG1659 	(WX11105,WX11104);
	dff 	XG1660 	(WX11107,WX11106);
	dff 	XG1661 	(WX11109,WX11108);
	dff 	XG1662 	(WX11111,WX11110);
	dff 	XG1663 	(WX11113,WX11112);
	dff 	XG1664 	(WX11115,WX11114);
	dff 	XG1665 	(WX11117,WX11116);
	dff 	XG1666 	(WX11119,WX11118);
	dff 	XG1667 	(WX11121,WX11120);
	dff 	XG1668 	(WX11123,WX11122);
	dff 	XG1669 	(WX11125,WX11124);
	dff 	XG1670 	(WX11127,WX11126);
	dff 	XG1671 	(WX11129,WX11128);
	dff 	XG1672 	(WX11131,WX11130);
	dff 	XG1673 	(WX11133,WX11132);
	dff 	XG1674 	(WX11135,WX11134);
	dff 	XG1675 	(WX11137,WX11136);
	dff 	XG1676 	(WX11139,WX11138);
	dff 	XG1677 	(WX11141,WX11140);
	dff 	XG1678 	(WX11143,WX11142);
	dff 	XG1679 	(WX11145,WX11144);
	dff 	XG1680 	(WX11147,WX11146);
	dff 	XG1681 	(WX11149,WX11148);
	dff 	XG1682 	(WX11151,WX11150);
	dff 	XG1683 	(WX11153,WX11152);
	dff 	XG1684 	(WX11155,WX11154);
	dff 	XG1685 	(WX11157,WX11156);
	dff 	XG1686 	(WX11159,WX11158);
	dff 	XG1687 	(WX11161,WX11160);
	dff 	XG1688 	(WX11163,WX11162);
	dff 	XG1689 	(WX11165,WX11164);
	dff 	XG1690 	(WX11167,WX11166);
	dff 	XG1691 	(WX11169,WX11168);
	dff 	XG1692 	(WX11171,WX11170);
	dff 	XG1693 	(WX11173,WX11172);
	dff 	XG1694 	(WX11175,WX11174);
	dff 	XG1695 	(WX11177,WX11176);
	dff 	XG1696 	(WX11179,WX11178);
	dff 	XG1697 	(WX11181,WX11180);
	dff 	XG1698 	(WX11183,WX11182);
	dff 	XG1699 	(WX11185,WX11184);
	dff 	XG1700 	(WX11187,WX11186);
	dff 	XG1701 	(WX11189,WX11188);
	dff 	XG1702 	(WX11191,WX11190);
	dff 	XG1703 	(WX11193,WX11192);
	dff 	XG1704 	(WX11195,WX11194);
	dff 	XG1705 	(WX11197,WX11196);
	dff 	XG1706 	(WX11199,WX11198);
	dff 	XG1707 	(WX11201,WX11200);
	dff 	XG1708 	(WX11203,WX11202);
	dff 	XG1709 	(WX11205,WX11204);
	dff 	XG1710 	(WX11207,WX11206);
	dff 	XG1711 	(WX11209,WX11208);
	dff 	XG1712 	(WX11211,WX11210);
	dff 	XG1713 	(WX11213,WX11212);
	dff 	XG1714 	(WX11215,WX11214);
	dff 	XG1715 	(WX11217,WX11216);
	dff 	XG1716 	(WX11219,WX11218);
	dff 	XG1717 	(WX11221,WX11220);
	dff 	XG1718 	(WX11223,WX11222);
	dff 	XG1719 	(WX11225,WX11224);
	dff 	XG1720 	(WX11227,WX11226);
	dff 	XG1721 	(WX11229,WX11228);
	dff 	XG1722 	(WX11231,WX11230);
	dff 	XG1723 	(WX11233,WX11232);
	dff 	XG1724 	(WX11235,WX11234);
	dff 	XG1725 	(WX11237,WX11236);
	dff 	XG1726 	(WX11239,WX11238);
	dff 	XG1727 	(WX11241,WX11240);
	dff 	XG1728 	(WX11243,WX11242);
	not 	XG1729 	(WX11574,RESET);
	not 	XG1730 	(WX10281,RESET);
	not 	XG1731 	(WX8988,RESET);
	not 	XG1732 	(WX7695,RESET);
	not 	XG1733 	(WX6402,RESET);
	not 	XG1734 	(WX5109,RESET);
	not 	XG1735 	(WX3816,RESET);
	not 	XG1736 	(WX2523,RESET);
	not 	XG1737 	(WX1230,RESET);
	not 	XG1738 	(WX11344,TM1);
	not 	XG1739 	(WX11343,TM1);
	not 	XG1740 	(WX10051,TM1);
	not 	XG1741 	(WX10050,TM1);
	not 	XG1742 	(WX8758,TM1);
	not 	XG1743 	(WX8757,TM1);
	not 	XG1744 	(WX7465,TM1);
	not 	XG1745 	(WX7464,TM1);
	not 	XG1746 	(WX6172,TM1);
	not 	XG1747 	(WX6171,TM1);
	not 	XG1748 	(WX4879,TM1);
	not 	XG1749 	(WX4878,TM1);
	not 	XG1750 	(WX3586,TM1);
	not 	XG1751 	(WX3585,TM1);
	not 	XG1752 	(WX2293,TM1);
	not 	XG1753 	(WX2292,TM1);
	not 	XG1754 	(WX1000,TM1);
	not 	XG1755 	(WX999,TM1);
	not 	XG1756 	(WX11342,TM0);
	not 	XG1757 	(WX11341,TM0);
	not 	XG1758 	(WX11340,TM0);
	not 	XG1759 	(WX10049,TM0);
	not 	XG1760 	(WX10048,TM0);
	not 	XG1761 	(WX10047,TM0);
	not 	XG1762 	(WX8756,TM0);
	not 	XG1763 	(WX8755,TM0);
	not 	XG1764 	(WX8754,TM0);
	not 	XG1765 	(WX7463,TM0);
	not 	XG1766 	(WX7462,TM0);
	not 	XG1767 	(WX7461,TM0);
	not 	XG1768 	(WX6170,TM0);
	not 	XG1769 	(WX6169,TM0);
	not 	XG1770 	(WX6168,TM0);
	not 	XG1771 	(WX4877,TM0);
	not 	XG1772 	(WX4876,TM0);
	not 	XG1773 	(WX4875,TM0);
	not 	XG1774 	(WX3584,TM0);
	not 	XG1775 	(WX3583,TM0);
	not 	XG1776 	(WX3582,TM0);
	not 	XG1777 	(WX2291,TM0);
	not 	XG1778 	(WX2290,TM0);
	not 	XG1779 	(WX2289,TM0);
	not 	XG1780 	(WX998,TM0);
	not 	XG1781 	(WX997,TM0);
	not 	XG1782 	(WX996,TM0);
	not 	XG1783 	(WX1005,WX996);
	not 	XG1784 	(WX1004,WX997);
	not 	XG1785 	(WX1002,WX998);
	not 	XG1786 	(WX2298,WX2289);
	not 	XG1787 	(WX2297,WX2290);
	not 	XG1788 	(WX2295,WX2291);
	not 	XG1789 	(WX3591,WX3582);
	not 	XG1790 	(WX3590,WX3583);
	not 	XG1791 	(WX3588,WX3584);
	not 	XG1792 	(WX4884,WX4875);
	not 	XG1793 	(WX4883,WX4876);
	not 	XG1794 	(WX4881,WX4877);
	not 	XG1795 	(WX6177,WX6168);
	not 	XG1796 	(WX6176,WX6169);
	not 	XG1797 	(WX6174,WX6170);
	not 	XG1798 	(WX7470,WX7461);
	not 	XG1799 	(WX7469,WX7462);
	not 	XG1800 	(WX7467,WX7463);
	not 	XG1801 	(WX8763,WX8754);
	not 	XG1802 	(WX8762,WX8755);
	not 	XG1803 	(WX8760,WX8756);
	not 	XG1804 	(WX10056,WX10047);
	not 	XG1805 	(WX10055,WX10048);
	not 	XG1806 	(WX10053,WX10049);
	not 	XG1807 	(WX11349,WX11340);
	not 	XG1808 	(WX11348,WX11341);
	not 	XG1809 	(WX11346,WX11342);
	not 	XG1810 	(WX1003,WX999);
	not 	XG1811 	(WX1001,WX1000);
	not 	XG1812 	(WX2296,WX2292);
	not 	XG1813 	(WX2294,WX2293);
	not 	XG1814 	(WX3589,WX3585);
	not 	XG1815 	(WX3587,WX3586);
	not 	XG1816 	(WX4882,WX4878);
	not 	XG1817 	(WX4880,WX4879);
	not 	XG1818 	(WX6175,WX6171);
	not 	XG1819 	(WX6173,WX6172);
	not 	XG1820 	(WX7468,WX7464);
	not 	XG1821 	(WX7466,WX7465);
	not 	XG1822 	(WX8761,WX8757);
	not 	XG1823 	(WX8759,WX8758);
	not 	XG1824 	(WX10054,WX10050);
	not 	XG1825 	(WX10052,WX10051);
	not 	XG1826 	(WX11347,WX11343);
	not 	XG1827 	(WX11345,WX11344);
	not 	XG1828 	(WX1263,WX1230);
	not 	XG1829 	(WX2556,WX2523);
	not 	XG1830 	(WX3849,WX3816);
	not 	XG1831 	(WX5142,WX5109);
	not 	XG1832 	(WX6435,WX6402);
	not 	XG1833 	(WX7728,WX7695);
	not 	XG1834 	(WX9021,WX8988);
	not 	XG1835 	(WX10314,WX10281);
	not 	XG1836 	(WX11607,WX11574);
	and 	XG1837 	(WX11242,RESET,WX11179);
	and 	XG1838 	(WX11240,RESET,WX11177);
	and 	XG1839 	(WX11238,RESET,WX11175);
	and 	XG1840 	(WX11236,RESET,WX11173);
	and 	XG1841 	(WX11234,RESET,WX11171);
	and 	XG1842 	(WX11232,RESET,WX11169);
	and 	XG1843 	(WX11230,RESET,WX11167);
	and 	XG1844 	(WX11228,RESET,WX11165);
	and 	XG1845 	(WX11226,RESET,WX11163);
	and 	XG1846 	(WX11224,RESET,WX11161);
	and 	XG1847 	(WX11222,RESET,WX11159);
	and 	XG1848 	(WX11220,RESET,WX11157);
	and 	XG1849 	(WX11218,RESET,WX11155);
	and 	XG1850 	(WX11216,RESET,WX11153);
	and 	XG1851 	(WX11214,RESET,WX11151);
	and 	XG1852 	(WX11212,RESET,WX11149);
	and 	XG1853 	(WX11210,RESET,WX11147);
	and 	XG1854 	(WX11208,RESET,WX11145);
	and 	XG1855 	(WX11206,RESET,WX11143);
	and 	XG1856 	(WX11204,RESET,WX11141);
	and 	XG1857 	(WX11202,RESET,WX11139);
	and 	XG1858 	(WX11200,RESET,WX11137);
	and 	XG1859 	(WX11198,RESET,WX11135);
	and 	XG1860 	(WX11196,RESET,WX11133);
	and 	XG1861 	(WX11194,RESET,WX11131);
	and 	XG1862 	(WX11192,RESET,WX11129);
	and 	XG1863 	(WX11190,RESET,WX11127);
	and 	XG1864 	(WX11188,RESET,WX11125);
	and 	XG1865 	(WX11186,RESET,WX11123);
	and 	XG1866 	(WX11184,RESET,WX11121);
	and 	XG1867 	(WX11182,RESET,WX11119);
	and 	XG1868 	(WX11180,RESET,WX11117);
	and 	XG1869 	(WX11178,RESET,WX11115);
	and 	XG1870 	(WX11176,RESET,WX11113);
	and 	XG1871 	(WX11174,RESET,WX11111);
	and 	XG1872 	(WX11172,RESET,WX11109);
	and 	XG1873 	(WX11170,RESET,WX11107);
	and 	XG1874 	(WX11168,RESET,WX11105);
	and 	XG1875 	(WX11166,RESET,WX11103);
	and 	XG1876 	(WX11164,RESET,WX11101);
	and 	XG1877 	(WX11162,RESET,WX11099);
	and 	XG1878 	(WX11160,RESET,WX11097);
	and 	XG1879 	(WX11158,RESET,WX11095);
	and 	XG1880 	(WX11156,RESET,WX11093);
	and 	XG1881 	(WX11154,RESET,WX11091);
	and 	XG1882 	(WX11152,RESET,WX11089);
	and 	XG1883 	(WX11150,RESET,WX11087);
	and 	XG1884 	(WX11148,RESET,WX11085);
	and 	XG1885 	(WX11146,RESET,WX11083);
	and 	XG1886 	(WX11144,RESET,WX11081);
	and 	XG1887 	(WX11142,RESET,WX11079);
	and 	XG1888 	(WX11140,RESET,WX11077);
	and 	XG1889 	(WX11138,RESET,WX11075);
	and 	XG1890 	(WX11136,RESET,WX11073);
	and 	XG1891 	(WX11134,RESET,WX11071);
	and 	XG1892 	(WX11132,RESET,WX11069);
	and 	XG1893 	(WX11130,RESET,WX11067);
	and 	XG1894 	(WX11128,RESET,WX11065);
	and 	XG1895 	(WX11126,RESET,WX11063);
	and 	XG1896 	(WX11124,RESET,WX11061);
	and 	XG1897 	(WX11122,RESET,WX11059);
	and 	XG1898 	(WX11120,RESET,WX11057);
	and 	XG1899 	(WX11118,RESET,WX11055);
	and 	XG1900 	(WX11116,RESET,WX11053);
	and 	XG1901 	(WX11114,RESET,WX11051);
	and 	XG1902 	(WX11112,RESET,WX11049);
	and 	XG1903 	(WX11110,RESET,WX11047);
	and 	XG1904 	(WX11108,RESET,WX11045);
	and 	XG1905 	(WX11106,RESET,WX11043);
	and 	XG1906 	(WX11104,RESET,WX11041);
	and 	XG1907 	(WX11102,RESET,WX11039);
	and 	XG1908 	(WX11100,RESET,WX11037);
	and 	XG1909 	(WX11098,RESET,WX11035);
	and 	XG1910 	(WX11096,RESET,WX11033);
	and 	XG1911 	(WX11094,RESET,WX11031);
	and 	XG1912 	(WX11092,RESET,WX11029);
	and 	XG1913 	(WX11090,RESET,WX11027);
	and 	XG1914 	(WX11088,RESET,WX11025);
	and 	XG1915 	(WX11086,RESET,WX11023);
	and 	XG1916 	(WX11084,RESET,WX11021);
	and 	XG1917 	(WX11082,RESET,WX11019);
	and 	XG1918 	(WX11080,RESET,WX11017);
	and 	XG1919 	(WX11078,RESET,WX11015);
	and 	XG1920 	(WX11076,RESET,WX11013);
	and 	XG1921 	(WX11074,RESET,WX11011);
	and 	XG1922 	(WX11072,RESET,WX11009);
	and 	XG1923 	(WX11070,RESET,WX11007);
	and 	XG1924 	(WX11068,RESET,WX11005);
	and 	XG1925 	(WX11066,RESET,WX11003);
	and 	XG1926 	(WX11064,RESET,WX11001);
	and 	XG1927 	(WX11062,RESET,WX10999);
	and 	XG1928 	(WX11060,RESET,WX10997);
	and 	XG1929 	(WX11058,RESET,WX10995);
	and 	XG1930 	(WX11056,RESET,WX10993);
	and 	XG1931 	(WX11054,RESET,WX10991);
	and 	XG1932 	(WX11052,RESET,WX10989);
	and 	XG1933 	(WX10888,RESET,WX10891);
	and 	XG1934 	(WX10886,RESET,WX10889);
	and 	XG1935 	(WX10884,RESET,WX10887);
	and 	XG1936 	(WX10882,RESET,WX10885);
	and 	XG1937 	(WX10880,RESET,WX10883);
	and 	XG1938 	(WX10878,RESET,WX10881);
	and 	XG1939 	(WX10876,RESET,WX10879);
	and 	XG1940 	(WX10874,RESET,WX10877);
	and 	XG1941 	(WX10872,RESET,WX10875);
	and 	XG1942 	(WX10870,RESET,WX10873);
	and 	XG1943 	(WX10868,RESET,WX10871);
	and 	XG1944 	(WX10866,RESET,WX10869);
	and 	XG1945 	(WX10864,RESET,WX10867);
	and 	XG1946 	(WX10862,RESET,WX10865);
	and 	XG1947 	(WX10860,RESET,WX10863);
	and 	XG1948 	(WX10858,RESET,WX10861);
	and 	XG1949 	(WX10856,RESET,WX10859);
	and 	XG1950 	(WX10854,RESET,WX10857);
	and 	XG1951 	(WX10852,RESET,WX10855);
	and 	XG1952 	(WX10850,RESET,WX10853);
	and 	XG1953 	(WX10848,RESET,WX10851);
	and 	XG1954 	(WX10846,RESET,WX10849);
	and 	XG1955 	(WX10844,RESET,WX10847);
	and 	XG1956 	(WX10842,RESET,WX10845);
	and 	XG1957 	(WX10840,RESET,WX10843);
	and 	XG1958 	(WX10838,RESET,WX10841);
	and 	XG1959 	(WX10836,RESET,WX10839);
	and 	XG1960 	(WX10834,RESET,WX10837);
	and 	XG1961 	(WX10832,RESET,WX10835);
	and 	XG1962 	(WX10830,RESET,WX10833);
	and 	XG1963 	(WX10828,RESET,WX10831);
	and 	XG1964 	(WX9949,RESET,WX9886);
	and 	XG1965 	(WX9947,RESET,WX9884);
	and 	XG1966 	(WX9945,RESET,WX9882);
	and 	XG1967 	(WX9943,RESET,WX9880);
	and 	XG1968 	(WX9941,RESET,WX9878);
	and 	XG1969 	(WX9939,RESET,WX9876);
	and 	XG1970 	(WX9937,RESET,WX9874);
	and 	XG1971 	(WX9935,RESET,WX9872);
	and 	XG1972 	(WX9933,RESET,WX9870);
	and 	XG1973 	(WX9931,RESET,WX9868);
	and 	XG1974 	(WX9929,RESET,WX9866);
	and 	XG1975 	(WX9927,RESET,WX9864);
	and 	XG1976 	(WX9925,RESET,WX9862);
	and 	XG1977 	(WX9923,RESET,WX9860);
	and 	XG1978 	(WX9921,RESET,WX9858);
	and 	XG1979 	(WX9919,RESET,WX9856);
	and 	XG1980 	(WX9917,RESET,WX9854);
	and 	XG1981 	(WX9915,RESET,WX9852);
	and 	XG1982 	(WX9913,RESET,WX9850);
	and 	XG1983 	(WX9911,RESET,WX9848);
	and 	XG1984 	(WX9909,RESET,WX9846);
	and 	XG1985 	(WX9907,RESET,WX9844);
	and 	XG1986 	(WX9905,RESET,WX9842);
	and 	XG1987 	(WX9903,RESET,WX9840);
	and 	XG1988 	(WX9901,RESET,WX9838);
	and 	XG1989 	(WX9899,RESET,WX9836);
	and 	XG1990 	(WX9897,RESET,WX9834);
	and 	XG1991 	(WX9895,RESET,WX9832);
	and 	XG1992 	(WX9893,RESET,WX9830);
	and 	XG1993 	(WX9891,RESET,WX9828);
	and 	XG1994 	(WX9889,RESET,WX9826);
	and 	XG1995 	(WX9887,RESET,WX9824);
	and 	XG1996 	(WX9885,RESET,WX9822);
	and 	XG1997 	(WX9883,RESET,WX9820);
	and 	XG1998 	(WX9881,RESET,WX9818);
	and 	XG1999 	(WX9879,RESET,WX9816);
	and 	XG2000 	(WX9877,RESET,WX9814);
	and 	XG2001 	(WX9875,RESET,WX9812);
	and 	XG2002 	(WX9873,RESET,WX9810);
	and 	XG2003 	(WX9871,RESET,WX9808);
	and 	XG2004 	(WX9869,RESET,WX9806);
	and 	XG2005 	(WX9867,RESET,WX9804);
	and 	XG2006 	(WX9865,RESET,WX9802);
	and 	XG2007 	(WX9863,RESET,WX9800);
	and 	XG2008 	(WX9861,RESET,WX9798);
	and 	XG2009 	(WX9859,RESET,WX9796);
	and 	XG2010 	(WX9857,RESET,WX9794);
	and 	XG2011 	(WX9855,RESET,WX9792);
	and 	XG2012 	(WX9853,RESET,WX9790);
	and 	XG2013 	(WX9851,RESET,WX9788);
	and 	XG2014 	(WX9849,RESET,WX9786);
	and 	XG2015 	(WX9847,RESET,WX9784);
	and 	XG2016 	(WX9845,RESET,WX9782);
	and 	XG2017 	(WX9843,RESET,WX9780);
	and 	XG2018 	(WX9841,RESET,WX9778);
	and 	XG2019 	(WX9839,RESET,WX9776);
	and 	XG2020 	(WX9837,RESET,WX9774);
	and 	XG2021 	(WX9835,RESET,WX9772);
	and 	XG2022 	(WX9833,RESET,WX9770);
	and 	XG2023 	(WX9831,RESET,WX9768);
	and 	XG2024 	(WX9829,RESET,WX9766);
	and 	XG2025 	(WX9827,RESET,WX9764);
	and 	XG2026 	(WX9825,RESET,WX9762);
	and 	XG2027 	(WX9823,RESET,WX9760);
	and 	XG2028 	(WX9821,RESET,WX9758);
	and 	XG2029 	(WX9819,RESET,WX9756);
	and 	XG2030 	(WX9817,RESET,WX9754);
	and 	XG2031 	(WX9815,RESET,WX9752);
	and 	XG2032 	(WX9813,RESET,WX9750);
	and 	XG2033 	(WX9811,RESET,WX9748);
	and 	XG2034 	(WX9809,RESET,WX9746);
	and 	XG2035 	(WX9807,RESET,WX9744);
	and 	XG2036 	(WX9805,RESET,WX9742);
	and 	XG2037 	(WX9803,RESET,WX9740);
	and 	XG2038 	(WX9801,RESET,WX9738);
	and 	XG2039 	(WX9799,RESET,WX9736);
	and 	XG2040 	(WX9797,RESET,WX9734);
	and 	XG2041 	(WX9795,RESET,WX9732);
	and 	XG2042 	(WX9793,RESET,WX9730);
	and 	XG2043 	(WX9791,RESET,WX9728);
	and 	XG2044 	(WX9789,RESET,WX9726);
	and 	XG2045 	(WX9787,RESET,WX9724);
	and 	XG2046 	(WX9785,RESET,WX9722);
	and 	XG2047 	(WX9783,RESET,WX9720);
	and 	XG2048 	(WX9781,RESET,WX9718);
	and 	XG2049 	(WX9779,RESET,WX9716);
	and 	XG2050 	(WX9777,RESET,WX9714);
	and 	XG2051 	(WX9775,RESET,WX9712);
	and 	XG2052 	(WX9773,RESET,WX9710);
	and 	XG2053 	(WX9771,RESET,WX9708);
	and 	XG2054 	(WX9769,RESET,WX9706);
	and 	XG2055 	(WX9767,RESET,WX9704);
	and 	XG2056 	(WX9765,RESET,WX9702);
	and 	XG2057 	(WX9763,RESET,WX9700);
	and 	XG2058 	(WX9761,RESET,WX9698);
	and 	XG2059 	(WX9759,RESET,WX9696);
	and 	XG2060 	(WX9595,RESET,WX9598);
	and 	XG2061 	(WX9593,RESET,WX9596);
	and 	XG2062 	(WX9591,RESET,WX9594);
	and 	XG2063 	(WX9589,RESET,WX9592);
	and 	XG2064 	(WX9587,RESET,WX9590);
	and 	XG2065 	(WX9585,RESET,WX9588);
	and 	XG2066 	(WX9583,RESET,WX9586);
	and 	XG2067 	(WX9581,RESET,WX9584);
	and 	XG2068 	(WX9579,RESET,WX9582);
	and 	XG2069 	(WX9577,RESET,WX9580);
	and 	XG2070 	(WX9575,RESET,WX9578);
	and 	XG2071 	(WX9573,RESET,WX9576);
	and 	XG2072 	(WX9571,RESET,WX9574);
	and 	XG2073 	(WX9569,RESET,WX9572);
	and 	XG2074 	(WX9567,RESET,WX9570);
	and 	XG2075 	(WX9565,RESET,WX9568);
	and 	XG2076 	(WX9563,RESET,WX9566);
	and 	XG2077 	(WX9561,RESET,WX9564);
	and 	XG2078 	(WX9559,RESET,WX9562);
	and 	XG2079 	(WX9557,RESET,WX9560);
	and 	XG2080 	(WX9555,RESET,WX9558);
	and 	XG2081 	(WX9553,RESET,WX9556);
	and 	XG2082 	(WX9551,RESET,WX9554);
	and 	XG2083 	(WX9549,RESET,WX9552);
	and 	XG2084 	(WX9547,RESET,WX9550);
	and 	XG2085 	(WX9545,RESET,WX9548);
	and 	XG2086 	(WX9543,RESET,WX9546);
	and 	XG2087 	(WX9541,RESET,WX9544);
	and 	XG2088 	(WX9539,RESET,WX9542);
	and 	XG2089 	(WX9537,RESET,WX9540);
	and 	XG2090 	(WX9535,RESET,WX9538);
	and 	XG2091 	(WX8656,RESET,WX8593);
	and 	XG2092 	(WX8654,RESET,WX8591);
	and 	XG2093 	(WX8652,RESET,WX8589);
	and 	XG2094 	(WX8650,RESET,WX8587);
	and 	XG2095 	(WX8648,RESET,WX8585);
	and 	XG2096 	(WX8646,RESET,WX8583);
	and 	XG2097 	(WX8644,RESET,WX8581);
	and 	XG2098 	(WX8642,RESET,WX8579);
	and 	XG2099 	(WX8640,RESET,WX8577);
	and 	XG2100 	(WX8638,RESET,WX8575);
	and 	XG2101 	(WX8636,RESET,WX8573);
	and 	XG2102 	(WX8634,RESET,WX8571);
	and 	XG2103 	(WX8632,RESET,WX8569);
	and 	XG2104 	(WX8630,RESET,WX8567);
	and 	XG2105 	(WX8628,RESET,WX8565);
	and 	XG2106 	(WX8626,RESET,WX8563);
	and 	XG2107 	(WX8624,RESET,WX8561);
	and 	XG2108 	(WX8622,RESET,WX8559);
	and 	XG2109 	(WX8620,RESET,WX8557);
	and 	XG2110 	(WX8618,RESET,WX8555);
	and 	XG2111 	(WX8616,RESET,WX8553);
	and 	XG2112 	(WX8614,RESET,WX8551);
	and 	XG2113 	(WX8612,RESET,WX8549);
	and 	XG2114 	(WX8610,RESET,WX8547);
	and 	XG2115 	(WX8608,RESET,WX8545);
	and 	XG2116 	(WX8606,RESET,WX8543);
	and 	XG2117 	(WX8604,RESET,WX8541);
	and 	XG2118 	(WX8602,RESET,WX8539);
	and 	XG2119 	(WX8600,RESET,WX8537);
	and 	XG2120 	(WX8598,RESET,WX8535);
	and 	XG2121 	(WX8596,RESET,WX8533);
	and 	XG2122 	(WX8594,RESET,WX8531);
	and 	XG2123 	(WX8592,RESET,WX8529);
	and 	XG2124 	(WX8590,RESET,WX8527);
	and 	XG2125 	(WX8588,RESET,WX8525);
	and 	XG2126 	(WX8586,RESET,WX8523);
	and 	XG2127 	(WX8584,RESET,WX8521);
	and 	XG2128 	(WX8582,RESET,WX8519);
	and 	XG2129 	(WX8580,RESET,WX8517);
	and 	XG2130 	(WX8578,RESET,WX8515);
	and 	XG2131 	(WX8576,RESET,WX8513);
	and 	XG2132 	(WX8574,RESET,WX8511);
	and 	XG2133 	(WX8572,RESET,WX8509);
	and 	XG2134 	(WX8570,RESET,WX8507);
	and 	XG2135 	(WX8568,RESET,WX8505);
	and 	XG2136 	(WX8566,RESET,WX8503);
	and 	XG2137 	(WX8564,RESET,WX8501);
	and 	XG2138 	(WX8562,RESET,WX8499);
	and 	XG2139 	(WX8560,RESET,WX8497);
	and 	XG2140 	(WX8558,RESET,WX8495);
	and 	XG2141 	(WX8556,RESET,WX8493);
	and 	XG2142 	(WX8554,RESET,WX8491);
	and 	XG2143 	(WX8552,RESET,WX8489);
	and 	XG2144 	(WX8550,RESET,WX8487);
	and 	XG2145 	(WX8548,RESET,WX8485);
	and 	XG2146 	(WX8546,RESET,WX8483);
	and 	XG2147 	(WX8544,RESET,WX8481);
	and 	XG2148 	(WX8542,RESET,WX8479);
	and 	XG2149 	(WX8540,RESET,WX8477);
	and 	XG2150 	(WX8538,RESET,WX8475);
	and 	XG2151 	(WX8536,RESET,WX8473);
	and 	XG2152 	(WX8534,RESET,WX8471);
	and 	XG2153 	(WX8532,RESET,WX8469);
	and 	XG2154 	(WX8530,RESET,WX8467);
	and 	XG2155 	(WX8528,RESET,WX8465);
	and 	XG2156 	(WX8526,RESET,WX8463);
	and 	XG2157 	(WX8524,RESET,WX8461);
	and 	XG2158 	(WX8522,RESET,WX8459);
	and 	XG2159 	(WX8520,RESET,WX8457);
	and 	XG2160 	(WX8518,RESET,WX8455);
	and 	XG2161 	(WX8516,RESET,WX8453);
	and 	XG2162 	(WX8514,RESET,WX8451);
	and 	XG2163 	(WX8512,RESET,WX8449);
	and 	XG2164 	(WX8510,RESET,WX8447);
	and 	XG2165 	(WX8508,RESET,WX8445);
	and 	XG2166 	(WX8506,RESET,WX8443);
	and 	XG2167 	(WX8504,RESET,WX8441);
	and 	XG2168 	(WX8502,RESET,WX8439);
	and 	XG2169 	(WX8500,RESET,WX8437);
	and 	XG2170 	(WX8498,RESET,WX8435);
	and 	XG2171 	(WX8496,RESET,WX8433);
	and 	XG2172 	(WX8494,RESET,WX8431);
	and 	XG2173 	(WX8492,RESET,WX8429);
	and 	XG2174 	(WX8490,RESET,WX8427);
	and 	XG2175 	(WX8488,RESET,WX8425);
	and 	XG2176 	(WX8486,RESET,WX8423);
	and 	XG2177 	(WX8484,RESET,WX8421);
	and 	XG2178 	(WX8482,RESET,WX8419);
	and 	XG2179 	(WX8480,RESET,WX8417);
	and 	XG2180 	(WX8478,RESET,WX8415);
	and 	XG2181 	(WX8476,RESET,WX8413);
	and 	XG2182 	(WX8474,RESET,WX8411);
	and 	XG2183 	(WX8472,RESET,WX8409);
	and 	XG2184 	(WX8470,RESET,WX8407);
	and 	XG2185 	(WX8468,RESET,WX8405);
	and 	XG2186 	(WX8466,RESET,WX8403);
	and 	XG2187 	(WX8302,RESET,WX8305);
	and 	XG2188 	(WX8300,RESET,WX8303);
	and 	XG2189 	(WX8298,RESET,WX8301);
	and 	XG2190 	(WX8296,RESET,WX8299);
	and 	XG2191 	(WX8294,RESET,WX8297);
	and 	XG2192 	(WX8292,RESET,WX8295);
	and 	XG2193 	(WX8290,RESET,WX8293);
	and 	XG2194 	(WX8288,RESET,WX8291);
	and 	XG2195 	(WX8286,RESET,WX8289);
	and 	XG2196 	(WX8284,RESET,WX8287);
	and 	XG2197 	(WX8282,RESET,WX8285);
	and 	XG2198 	(WX8280,RESET,WX8283);
	and 	XG2199 	(WX8278,RESET,WX8281);
	and 	XG2200 	(WX8276,RESET,WX8279);
	and 	XG2201 	(WX8274,RESET,WX8277);
	and 	XG2202 	(WX8272,RESET,WX8275);
	and 	XG2203 	(WX8270,RESET,WX8273);
	and 	XG2204 	(WX8268,RESET,WX8271);
	and 	XG2205 	(WX8266,RESET,WX8269);
	and 	XG2206 	(WX8264,RESET,WX8267);
	and 	XG2207 	(WX8262,RESET,WX8265);
	and 	XG2208 	(WX8260,RESET,WX8263);
	and 	XG2209 	(WX8258,RESET,WX8261);
	and 	XG2210 	(WX8256,RESET,WX8259);
	and 	XG2211 	(WX8254,RESET,WX8257);
	and 	XG2212 	(WX8252,RESET,WX8255);
	and 	XG2213 	(WX8250,RESET,WX8253);
	and 	XG2214 	(WX8248,RESET,WX8251);
	and 	XG2215 	(WX8246,RESET,WX8249);
	and 	XG2216 	(WX8244,RESET,WX8247);
	and 	XG2217 	(WX8242,RESET,WX8245);
	and 	XG2218 	(WX7363,RESET,WX7300);
	and 	XG2219 	(WX7361,RESET,WX7298);
	and 	XG2220 	(WX7359,RESET,WX7296);
	and 	XG2221 	(WX7357,RESET,WX7294);
	and 	XG2222 	(WX7355,RESET,WX7292);
	and 	XG2223 	(WX7353,RESET,WX7290);
	and 	XG2224 	(WX7351,RESET,WX7288);
	and 	XG2225 	(WX7349,RESET,WX7286);
	and 	XG2226 	(WX7347,RESET,WX7284);
	and 	XG2227 	(WX7345,RESET,WX7282);
	and 	XG2228 	(WX7343,RESET,WX7280);
	and 	XG2229 	(WX7341,RESET,WX7278);
	and 	XG2230 	(WX7339,RESET,WX7276);
	and 	XG2231 	(WX7337,RESET,WX7274);
	and 	XG2232 	(WX7335,RESET,WX7272);
	and 	XG2233 	(WX7333,RESET,WX7270);
	and 	XG2234 	(WX7331,RESET,WX7268);
	and 	XG2235 	(WX7329,RESET,WX7266);
	and 	XG2236 	(WX7327,RESET,WX7264);
	and 	XG2237 	(WX7325,RESET,WX7262);
	and 	XG2238 	(WX7323,RESET,WX7260);
	and 	XG2239 	(WX7321,RESET,WX7258);
	and 	XG2240 	(WX7319,RESET,WX7256);
	and 	XG2241 	(WX7317,RESET,WX7254);
	and 	XG2242 	(WX7315,RESET,WX7252);
	and 	XG2243 	(WX7313,RESET,WX7250);
	and 	XG2244 	(WX7311,RESET,WX7248);
	and 	XG2245 	(WX7309,RESET,WX7246);
	and 	XG2246 	(WX7307,RESET,WX7244);
	and 	XG2247 	(WX7305,RESET,WX7242);
	and 	XG2248 	(WX7303,RESET,WX7240);
	and 	XG2249 	(WX7301,RESET,WX7238);
	and 	XG2250 	(WX7299,RESET,WX7236);
	and 	XG2251 	(WX7297,RESET,WX7234);
	and 	XG2252 	(WX7295,RESET,WX7232);
	and 	XG2253 	(WX7293,RESET,WX7230);
	and 	XG2254 	(WX7291,RESET,WX7228);
	and 	XG2255 	(WX7289,RESET,WX7226);
	and 	XG2256 	(WX7287,RESET,WX7224);
	and 	XG2257 	(WX7285,RESET,WX7222);
	and 	XG2258 	(WX7283,RESET,WX7220);
	and 	XG2259 	(WX7281,RESET,WX7218);
	and 	XG2260 	(WX7279,RESET,WX7216);
	and 	XG2261 	(WX7277,RESET,WX7214);
	and 	XG2262 	(WX7275,RESET,WX7212);
	and 	XG2263 	(WX7273,RESET,WX7210);
	and 	XG2264 	(WX7271,RESET,WX7208);
	and 	XG2265 	(WX7269,RESET,WX7206);
	and 	XG2266 	(WX7267,RESET,WX7204);
	and 	XG2267 	(WX7265,RESET,WX7202);
	and 	XG2268 	(WX7263,RESET,WX7200);
	and 	XG2269 	(WX7261,RESET,WX7198);
	and 	XG2270 	(WX7259,RESET,WX7196);
	and 	XG2271 	(WX7257,RESET,WX7194);
	and 	XG2272 	(WX7255,RESET,WX7192);
	and 	XG2273 	(WX7253,RESET,WX7190);
	and 	XG2274 	(WX7251,RESET,WX7188);
	and 	XG2275 	(WX7249,RESET,WX7186);
	and 	XG2276 	(WX7247,RESET,WX7184);
	and 	XG2277 	(WX7245,RESET,WX7182);
	and 	XG2278 	(WX7243,RESET,WX7180);
	and 	XG2279 	(WX7241,RESET,WX7178);
	and 	XG2280 	(WX7239,RESET,WX7176);
	and 	XG2281 	(WX7237,RESET,WX7174);
	and 	XG2282 	(WX7235,RESET,WX7172);
	and 	XG2283 	(WX7233,RESET,WX7170);
	and 	XG2284 	(WX7231,RESET,WX7168);
	and 	XG2285 	(WX7229,RESET,WX7166);
	and 	XG2286 	(WX7227,RESET,WX7164);
	and 	XG2287 	(WX7225,RESET,WX7162);
	and 	XG2288 	(WX7223,RESET,WX7160);
	and 	XG2289 	(WX7221,RESET,WX7158);
	and 	XG2290 	(WX7219,RESET,WX7156);
	and 	XG2291 	(WX7217,RESET,WX7154);
	and 	XG2292 	(WX7215,RESET,WX7152);
	and 	XG2293 	(WX7213,RESET,WX7150);
	and 	XG2294 	(WX7211,RESET,WX7148);
	and 	XG2295 	(WX7209,RESET,WX7146);
	and 	XG2296 	(WX7207,RESET,WX7144);
	and 	XG2297 	(WX7205,RESET,WX7142);
	and 	XG2298 	(WX7203,RESET,WX7140);
	and 	XG2299 	(WX7201,RESET,WX7138);
	and 	XG2300 	(WX7199,RESET,WX7136);
	and 	XG2301 	(WX7197,RESET,WX7134);
	and 	XG2302 	(WX7195,RESET,WX7132);
	and 	XG2303 	(WX7193,RESET,WX7130);
	and 	XG2304 	(WX7191,RESET,WX7128);
	and 	XG2305 	(WX7189,RESET,WX7126);
	and 	XG2306 	(WX7187,RESET,WX7124);
	and 	XG2307 	(WX7185,RESET,WX7122);
	and 	XG2308 	(WX7183,RESET,WX7120);
	and 	XG2309 	(WX7181,RESET,WX7118);
	and 	XG2310 	(WX7179,RESET,WX7116);
	and 	XG2311 	(WX7177,RESET,WX7114);
	and 	XG2312 	(WX7175,RESET,WX7112);
	and 	XG2313 	(WX7173,RESET,WX7110);
	and 	XG2314 	(WX7009,RESET,WX7012);
	and 	XG2315 	(WX7007,RESET,WX7010);
	and 	XG2316 	(WX7005,RESET,WX7008);
	and 	XG2317 	(WX7003,RESET,WX7006);
	and 	XG2318 	(WX7001,RESET,WX7004);
	and 	XG2319 	(WX6999,RESET,WX7002);
	and 	XG2320 	(WX6997,RESET,WX7000);
	and 	XG2321 	(WX6995,RESET,WX6998);
	and 	XG2322 	(WX6993,RESET,WX6996);
	and 	XG2323 	(WX6991,RESET,WX6994);
	and 	XG2324 	(WX6989,RESET,WX6992);
	and 	XG2325 	(WX6987,RESET,WX6990);
	and 	XG2326 	(WX6985,RESET,WX6988);
	and 	XG2327 	(WX6983,RESET,WX6986);
	and 	XG2328 	(WX6981,RESET,WX6984);
	and 	XG2329 	(WX6979,RESET,WX6982);
	and 	XG2330 	(WX6977,RESET,WX6980);
	and 	XG2331 	(WX6975,RESET,WX6978);
	and 	XG2332 	(WX6973,RESET,WX6976);
	and 	XG2333 	(WX6971,RESET,WX6974);
	and 	XG2334 	(WX6969,RESET,WX6972);
	and 	XG2335 	(WX6967,RESET,WX6970);
	and 	XG2336 	(WX6965,RESET,WX6968);
	and 	XG2337 	(WX6963,RESET,WX6966);
	and 	XG2338 	(WX6961,RESET,WX6964);
	and 	XG2339 	(WX6959,RESET,WX6962);
	and 	XG2340 	(WX6957,RESET,WX6960);
	and 	XG2341 	(WX6955,RESET,WX6958);
	and 	XG2342 	(WX6953,RESET,WX6956);
	and 	XG2343 	(WX6951,RESET,WX6954);
	and 	XG2344 	(WX6949,RESET,WX6952);
	and 	XG2345 	(WX6070,RESET,WX6007);
	and 	XG2346 	(WX6068,RESET,WX6005);
	and 	XG2347 	(WX6066,RESET,WX6003);
	and 	XG2348 	(WX6064,RESET,WX6001);
	and 	XG2349 	(WX6062,RESET,WX5999);
	and 	XG2350 	(WX6060,RESET,WX5997);
	and 	XG2351 	(WX6058,RESET,WX5995);
	and 	XG2352 	(WX6056,RESET,WX5993);
	and 	XG2353 	(WX6054,RESET,WX5991);
	and 	XG2354 	(WX6052,RESET,WX5989);
	and 	XG2355 	(WX6050,RESET,WX5987);
	and 	XG2356 	(WX6048,RESET,WX5985);
	and 	XG2357 	(WX6046,RESET,WX5983);
	and 	XG2358 	(WX6044,RESET,WX5981);
	and 	XG2359 	(WX6042,RESET,WX5979);
	and 	XG2360 	(WX6040,RESET,WX5977);
	and 	XG2361 	(WX6038,RESET,WX5975);
	and 	XG2362 	(WX6036,RESET,WX5973);
	and 	XG2363 	(WX6034,RESET,WX5971);
	and 	XG2364 	(WX6032,RESET,WX5969);
	and 	XG2365 	(WX6030,RESET,WX5967);
	and 	XG2366 	(WX6028,RESET,WX5965);
	and 	XG2367 	(WX6026,RESET,WX5963);
	and 	XG2368 	(WX6024,RESET,WX5961);
	and 	XG2369 	(WX6022,RESET,WX5959);
	and 	XG2370 	(WX6020,RESET,WX5957);
	and 	XG2371 	(WX6018,RESET,WX5955);
	and 	XG2372 	(WX6016,RESET,WX5953);
	and 	XG2373 	(WX6014,RESET,WX5951);
	and 	XG2374 	(WX6012,RESET,WX5949);
	and 	XG2375 	(WX6010,RESET,WX5947);
	and 	XG2376 	(WX6008,RESET,WX5945);
	and 	XG2377 	(WX6006,RESET,WX5943);
	and 	XG2378 	(WX6004,RESET,WX5941);
	and 	XG2379 	(WX6002,RESET,WX5939);
	and 	XG2380 	(WX6000,RESET,WX5937);
	and 	XG2381 	(WX5998,RESET,WX5935);
	and 	XG2382 	(WX5996,RESET,WX5933);
	and 	XG2383 	(WX5994,RESET,WX5931);
	and 	XG2384 	(WX5992,RESET,WX5929);
	and 	XG2385 	(WX5990,RESET,WX5927);
	and 	XG2386 	(WX5988,RESET,WX5925);
	and 	XG2387 	(WX5986,RESET,WX5923);
	and 	XG2388 	(WX5984,RESET,WX5921);
	and 	XG2389 	(WX5982,RESET,WX5919);
	and 	XG2390 	(WX5980,RESET,WX5917);
	and 	XG2391 	(WX5978,RESET,WX5915);
	and 	XG2392 	(WX5976,RESET,WX5913);
	and 	XG2393 	(WX5974,RESET,WX5911);
	and 	XG2394 	(WX5972,RESET,WX5909);
	and 	XG2395 	(WX5970,RESET,WX5907);
	and 	XG2396 	(WX5968,RESET,WX5905);
	and 	XG2397 	(WX5966,RESET,WX5903);
	and 	XG2398 	(WX5964,RESET,WX5901);
	and 	XG2399 	(WX5962,RESET,WX5899);
	and 	XG2400 	(WX5960,RESET,WX5897);
	and 	XG2401 	(WX5958,RESET,WX5895);
	and 	XG2402 	(WX5956,RESET,WX5893);
	and 	XG2403 	(WX5954,RESET,WX5891);
	and 	XG2404 	(WX5952,RESET,WX5889);
	and 	XG2405 	(WX5950,RESET,WX5887);
	and 	XG2406 	(WX5948,RESET,WX5885);
	and 	XG2407 	(WX5946,RESET,WX5883);
	and 	XG2408 	(WX5944,RESET,WX5881);
	and 	XG2409 	(WX5942,RESET,WX5879);
	and 	XG2410 	(WX5940,RESET,WX5877);
	and 	XG2411 	(WX5938,RESET,WX5875);
	and 	XG2412 	(WX5936,RESET,WX5873);
	and 	XG2413 	(WX5934,RESET,WX5871);
	and 	XG2414 	(WX5932,RESET,WX5869);
	and 	XG2415 	(WX5930,RESET,WX5867);
	and 	XG2416 	(WX5928,RESET,WX5865);
	and 	XG2417 	(WX5926,RESET,WX5863);
	and 	XG2418 	(WX5924,RESET,WX5861);
	and 	XG2419 	(WX5922,RESET,WX5859);
	and 	XG2420 	(WX5920,RESET,WX5857);
	and 	XG2421 	(WX5918,RESET,WX5855);
	and 	XG2422 	(WX5916,RESET,WX5853);
	and 	XG2423 	(WX5914,RESET,WX5851);
	and 	XG2424 	(WX5912,RESET,WX5849);
	and 	XG2425 	(WX5910,RESET,WX5847);
	and 	XG2426 	(WX5908,RESET,WX5845);
	and 	XG2427 	(WX5906,RESET,WX5843);
	and 	XG2428 	(WX5904,RESET,WX5841);
	and 	XG2429 	(WX5902,RESET,WX5839);
	and 	XG2430 	(WX5900,RESET,WX5837);
	and 	XG2431 	(WX5898,RESET,WX5835);
	and 	XG2432 	(WX5896,RESET,WX5833);
	and 	XG2433 	(WX5894,RESET,WX5831);
	and 	XG2434 	(WX5892,RESET,WX5829);
	and 	XG2435 	(WX5890,RESET,WX5827);
	and 	XG2436 	(WX5888,RESET,WX5825);
	and 	XG2437 	(WX5886,RESET,WX5823);
	and 	XG2438 	(WX5884,RESET,WX5821);
	and 	XG2439 	(WX5882,RESET,WX5819);
	and 	XG2440 	(WX5880,RESET,WX5817);
	and 	XG2441 	(WX5716,RESET,WX5719);
	and 	XG2442 	(WX5714,RESET,WX5717);
	and 	XG2443 	(WX5712,RESET,WX5715);
	and 	XG2444 	(WX5710,RESET,WX5713);
	and 	XG2445 	(WX5708,RESET,WX5711);
	and 	XG2446 	(WX5706,RESET,WX5709);
	and 	XG2447 	(WX5704,RESET,WX5707);
	and 	XG2448 	(WX5702,RESET,WX5705);
	and 	XG2449 	(WX5700,RESET,WX5703);
	and 	XG2450 	(WX5698,RESET,WX5701);
	and 	XG2451 	(WX5696,RESET,WX5699);
	and 	XG2452 	(WX5694,RESET,WX5697);
	and 	XG2453 	(WX5692,RESET,WX5695);
	and 	XG2454 	(WX5690,RESET,WX5693);
	and 	XG2455 	(WX5688,RESET,WX5691);
	and 	XG2456 	(WX5686,RESET,WX5689);
	and 	XG2457 	(WX5684,RESET,WX5687);
	and 	XG2458 	(WX5682,RESET,WX5685);
	and 	XG2459 	(WX5680,RESET,WX5683);
	and 	XG2460 	(WX5678,RESET,WX5681);
	and 	XG2461 	(WX5676,RESET,WX5679);
	and 	XG2462 	(WX5674,RESET,WX5677);
	and 	XG2463 	(WX5672,RESET,WX5675);
	and 	XG2464 	(WX5670,RESET,WX5673);
	and 	XG2465 	(WX5668,RESET,WX5671);
	and 	XG2466 	(WX5666,RESET,WX5669);
	and 	XG2467 	(WX5664,RESET,WX5667);
	and 	XG2468 	(WX5662,RESET,WX5665);
	and 	XG2469 	(WX5660,RESET,WX5663);
	and 	XG2470 	(WX5658,RESET,WX5661);
	and 	XG2471 	(WX5656,RESET,WX5659);
	and 	XG2472 	(WX4777,RESET,WX4714);
	and 	XG2473 	(WX4775,RESET,WX4712);
	and 	XG2474 	(WX4773,RESET,WX4710);
	and 	XG2475 	(WX4771,RESET,WX4708);
	and 	XG2476 	(WX4769,RESET,WX4706);
	and 	XG2477 	(WX4767,RESET,WX4704);
	and 	XG2478 	(WX4765,RESET,WX4702);
	and 	XG2479 	(WX4763,RESET,WX4700);
	and 	XG2480 	(WX4761,RESET,WX4698);
	and 	XG2481 	(WX4759,RESET,WX4696);
	and 	XG2482 	(WX4757,RESET,WX4694);
	and 	XG2483 	(WX4755,RESET,WX4692);
	and 	XG2484 	(WX4753,RESET,WX4690);
	and 	XG2485 	(WX4751,RESET,WX4688);
	and 	XG2486 	(WX4749,RESET,WX4686);
	and 	XG2487 	(WX4747,RESET,WX4684);
	and 	XG2488 	(WX4745,RESET,WX4682);
	and 	XG2489 	(WX4743,RESET,WX4680);
	and 	XG2490 	(WX4741,RESET,WX4678);
	and 	XG2491 	(WX4739,RESET,WX4676);
	and 	XG2492 	(WX4737,RESET,WX4674);
	and 	XG2493 	(WX4735,RESET,WX4672);
	and 	XG2494 	(WX4733,RESET,WX4670);
	and 	XG2495 	(WX4731,RESET,WX4668);
	and 	XG2496 	(WX4729,RESET,WX4666);
	and 	XG2497 	(WX4727,RESET,WX4664);
	and 	XG2498 	(WX4725,RESET,WX4662);
	and 	XG2499 	(WX4723,RESET,WX4660);
	and 	XG2500 	(WX4721,RESET,WX4658);
	and 	XG2501 	(WX4719,RESET,WX4656);
	and 	XG2502 	(WX4717,RESET,WX4654);
	and 	XG2503 	(WX4715,RESET,WX4652);
	and 	XG2504 	(WX4713,RESET,WX4650);
	and 	XG2505 	(WX4711,RESET,WX4648);
	and 	XG2506 	(WX4709,RESET,WX4646);
	and 	XG2507 	(WX4707,RESET,WX4644);
	and 	XG2508 	(WX4705,RESET,WX4642);
	and 	XG2509 	(WX4703,RESET,WX4640);
	and 	XG2510 	(WX4701,RESET,WX4638);
	and 	XG2511 	(WX4699,RESET,WX4636);
	and 	XG2512 	(WX4697,RESET,WX4634);
	and 	XG2513 	(WX4695,RESET,WX4632);
	and 	XG2514 	(WX4693,RESET,WX4630);
	and 	XG2515 	(WX4691,RESET,WX4628);
	and 	XG2516 	(WX4689,RESET,WX4626);
	and 	XG2517 	(WX4687,RESET,WX4624);
	and 	XG2518 	(WX4685,RESET,WX4622);
	and 	XG2519 	(WX4683,RESET,WX4620);
	and 	XG2520 	(WX4681,RESET,WX4618);
	and 	XG2521 	(WX4679,RESET,WX4616);
	and 	XG2522 	(WX4677,RESET,WX4614);
	and 	XG2523 	(WX4675,RESET,WX4612);
	and 	XG2524 	(WX4673,RESET,WX4610);
	and 	XG2525 	(WX4671,RESET,WX4608);
	and 	XG2526 	(WX4669,RESET,WX4606);
	and 	XG2527 	(WX4667,RESET,WX4604);
	and 	XG2528 	(WX4665,RESET,WX4602);
	and 	XG2529 	(WX4663,RESET,WX4600);
	and 	XG2530 	(WX4661,RESET,WX4598);
	and 	XG2531 	(WX4659,RESET,WX4596);
	and 	XG2532 	(WX4657,RESET,WX4594);
	and 	XG2533 	(WX4655,RESET,WX4592);
	and 	XG2534 	(WX4653,RESET,WX4590);
	and 	XG2535 	(WX4651,RESET,WX4588);
	and 	XG2536 	(WX4649,RESET,WX4586);
	and 	XG2537 	(WX4647,RESET,WX4584);
	and 	XG2538 	(WX4645,RESET,WX4582);
	and 	XG2539 	(WX4643,RESET,WX4580);
	and 	XG2540 	(WX4641,RESET,WX4578);
	and 	XG2541 	(WX4639,RESET,WX4576);
	and 	XG2542 	(WX4637,RESET,WX4574);
	and 	XG2543 	(WX4635,RESET,WX4572);
	and 	XG2544 	(WX4633,RESET,WX4570);
	and 	XG2545 	(WX4631,RESET,WX4568);
	and 	XG2546 	(WX4629,RESET,WX4566);
	and 	XG2547 	(WX4627,RESET,WX4564);
	and 	XG2548 	(WX4625,RESET,WX4562);
	and 	XG2549 	(WX4623,RESET,WX4560);
	and 	XG2550 	(WX4621,RESET,WX4558);
	and 	XG2551 	(WX4619,RESET,WX4556);
	and 	XG2552 	(WX4617,RESET,WX4554);
	and 	XG2553 	(WX4615,RESET,WX4552);
	and 	XG2554 	(WX4613,RESET,WX4550);
	and 	XG2555 	(WX4611,RESET,WX4548);
	and 	XG2556 	(WX4609,RESET,WX4546);
	and 	XG2557 	(WX4607,RESET,WX4544);
	and 	XG2558 	(WX4605,RESET,WX4542);
	and 	XG2559 	(WX4603,RESET,WX4540);
	and 	XG2560 	(WX4601,RESET,WX4538);
	and 	XG2561 	(WX4599,RESET,WX4536);
	and 	XG2562 	(WX4597,RESET,WX4534);
	and 	XG2563 	(WX4595,RESET,WX4532);
	and 	XG2564 	(WX4593,RESET,WX4530);
	and 	XG2565 	(WX4591,RESET,WX4528);
	and 	XG2566 	(WX4589,RESET,WX4526);
	and 	XG2567 	(WX4587,RESET,WX4524);
	and 	XG2568 	(WX4423,RESET,WX4426);
	and 	XG2569 	(WX4421,RESET,WX4424);
	and 	XG2570 	(WX4419,RESET,WX4422);
	and 	XG2571 	(WX4417,RESET,WX4420);
	and 	XG2572 	(WX4415,RESET,WX4418);
	and 	XG2573 	(WX4413,RESET,WX4416);
	and 	XG2574 	(WX4411,RESET,WX4414);
	and 	XG2575 	(WX4409,RESET,WX4412);
	and 	XG2576 	(WX4407,RESET,WX4410);
	and 	XG2577 	(WX4405,RESET,WX4408);
	and 	XG2578 	(WX4403,RESET,WX4406);
	and 	XG2579 	(WX4401,RESET,WX4404);
	and 	XG2580 	(WX4399,RESET,WX4402);
	and 	XG2581 	(WX4397,RESET,WX4400);
	and 	XG2582 	(WX4395,RESET,WX4398);
	and 	XG2583 	(WX4393,RESET,WX4396);
	and 	XG2584 	(WX4391,RESET,WX4394);
	and 	XG2585 	(WX4389,RESET,WX4392);
	and 	XG2586 	(WX4387,RESET,WX4390);
	and 	XG2587 	(WX4385,RESET,WX4388);
	and 	XG2588 	(WX4383,RESET,WX4386);
	and 	XG2589 	(WX4381,RESET,WX4384);
	and 	XG2590 	(WX4379,RESET,WX4382);
	and 	XG2591 	(WX4377,RESET,WX4380);
	and 	XG2592 	(WX4375,RESET,WX4378);
	and 	XG2593 	(WX4373,RESET,WX4376);
	and 	XG2594 	(WX4371,RESET,WX4374);
	and 	XG2595 	(WX4369,RESET,WX4372);
	and 	XG2596 	(WX4367,RESET,WX4370);
	and 	XG2597 	(WX4365,RESET,WX4368);
	and 	XG2598 	(WX4363,RESET,WX4366);
	and 	XG2599 	(WX3484,RESET,WX3421);
	and 	XG2600 	(WX3482,RESET,WX3419);
	and 	XG2601 	(WX3480,RESET,WX3417);
	and 	XG2602 	(WX3478,RESET,WX3415);
	and 	XG2603 	(WX3476,RESET,WX3413);
	and 	XG2604 	(WX3474,RESET,WX3411);
	and 	XG2605 	(WX3472,RESET,WX3409);
	and 	XG2606 	(WX3470,RESET,WX3407);
	and 	XG2607 	(WX3468,RESET,WX3405);
	and 	XG2608 	(WX3466,RESET,WX3403);
	and 	XG2609 	(WX3464,RESET,WX3401);
	and 	XG2610 	(WX3462,RESET,WX3399);
	and 	XG2611 	(WX3460,RESET,WX3397);
	and 	XG2612 	(WX3458,RESET,WX3395);
	and 	XG2613 	(WX3456,RESET,WX3393);
	and 	XG2614 	(WX3454,RESET,WX3391);
	and 	XG2615 	(WX3452,RESET,WX3389);
	and 	XG2616 	(WX3450,RESET,WX3387);
	and 	XG2617 	(WX3448,RESET,WX3385);
	and 	XG2618 	(WX3446,RESET,WX3383);
	and 	XG2619 	(WX3444,RESET,WX3381);
	and 	XG2620 	(WX3442,RESET,WX3379);
	and 	XG2621 	(WX3440,RESET,WX3377);
	and 	XG2622 	(WX3438,RESET,WX3375);
	and 	XG2623 	(WX3436,RESET,WX3373);
	and 	XG2624 	(WX3434,RESET,WX3371);
	and 	XG2625 	(WX3432,RESET,WX3369);
	and 	XG2626 	(WX3430,RESET,WX3367);
	and 	XG2627 	(WX3428,RESET,WX3365);
	and 	XG2628 	(WX3426,RESET,WX3363);
	and 	XG2629 	(WX3424,RESET,WX3361);
	and 	XG2630 	(WX3422,RESET,WX3359);
	and 	XG2631 	(WX3420,RESET,WX3357);
	and 	XG2632 	(WX3418,RESET,WX3355);
	and 	XG2633 	(WX3416,RESET,WX3353);
	and 	XG2634 	(WX3414,RESET,WX3351);
	and 	XG2635 	(WX3412,RESET,WX3349);
	and 	XG2636 	(WX3410,RESET,WX3347);
	and 	XG2637 	(WX3408,RESET,WX3345);
	and 	XG2638 	(WX3406,RESET,WX3343);
	and 	XG2639 	(WX3404,RESET,WX3341);
	and 	XG2640 	(WX3402,RESET,WX3339);
	and 	XG2641 	(WX3400,RESET,WX3337);
	and 	XG2642 	(WX3398,RESET,WX3335);
	and 	XG2643 	(WX3396,RESET,WX3333);
	and 	XG2644 	(WX3394,RESET,WX3331);
	and 	XG2645 	(WX3392,RESET,WX3329);
	and 	XG2646 	(WX3390,RESET,WX3327);
	and 	XG2647 	(WX3388,RESET,WX3325);
	and 	XG2648 	(WX3386,RESET,WX3323);
	and 	XG2649 	(WX3384,RESET,WX3321);
	and 	XG2650 	(WX3382,RESET,WX3319);
	and 	XG2651 	(WX3380,RESET,WX3317);
	and 	XG2652 	(WX3378,RESET,WX3315);
	and 	XG2653 	(WX3376,RESET,WX3313);
	and 	XG2654 	(WX3374,RESET,WX3311);
	and 	XG2655 	(WX3372,RESET,WX3309);
	and 	XG2656 	(WX3370,RESET,WX3307);
	and 	XG2657 	(WX3368,RESET,WX3305);
	and 	XG2658 	(WX3366,RESET,WX3303);
	and 	XG2659 	(WX3364,RESET,WX3301);
	and 	XG2660 	(WX3362,RESET,WX3299);
	and 	XG2661 	(WX3360,RESET,WX3297);
	and 	XG2662 	(WX3358,RESET,WX3295);
	and 	XG2663 	(WX3356,RESET,WX3293);
	and 	XG2664 	(WX3354,RESET,WX3291);
	and 	XG2665 	(WX3352,RESET,WX3289);
	and 	XG2666 	(WX3350,RESET,WX3287);
	and 	XG2667 	(WX3348,RESET,WX3285);
	and 	XG2668 	(WX3346,RESET,WX3283);
	and 	XG2669 	(WX3344,RESET,WX3281);
	and 	XG2670 	(WX3342,RESET,WX3279);
	and 	XG2671 	(WX3340,RESET,WX3277);
	and 	XG2672 	(WX3338,RESET,WX3275);
	and 	XG2673 	(WX3336,RESET,WX3273);
	and 	XG2674 	(WX3334,RESET,WX3271);
	and 	XG2675 	(WX3332,RESET,WX3269);
	and 	XG2676 	(WX3330,RESET,WX3267);
	and 	XG2677 	(WX3328,RESET,WX3265);
	and 	XG2678 	(WX3326,RESET,WX3263);
	and 	XG2679 	(WX3324,RESET,WX3261);
	and 	XG2680 	(WX3322,RESET,WX3259);
	and 	XG2681 	(WX3320,RESET,WX3257);
	and 	XG2682 	(WX3318,RESET,WX3255);
	and 	XG2683 	(WX3316,RESET,WX3253);
	and 	XG2684 	(WX3314,RESET,WX3251);
	and 	XG2685 	(WX3312,RESET,WX3249);
	and 	XG2686 	(WX3310,RESET,WX3247);
	and 	XG2687 	(WX3308,RESET,WX3245);
	and 	XG2688 	(WX3306,RESET,WX3243);
	and 	XG2689 	(WX3304,RESET,WX3241);
	and 	XG2690 	(WX3302,RESET,WX3239);
	and 	XG2691 	(WX3300,RESET,WX3237);
	and 	XG2692 	(WX3298,RESET,WX3235);
	and 	XG2693 	(WX3296,RESET,WX3233);
	and 	XG2694 	(WX3294,RESET,WX3231);
	and 	XG2695 	(WX3130,RESET,WX3133);
	and 	XG2696 	(WX3128,RESET,WX3131);
	and 	XG2697 	(WX3126,RESET,WX3129);
	and 	XG2698 	(WX3124,RESET,WX3127);
	and 	XG2699 	(WX3122,RESET,WX3125);
	and 	XG2700 	(WX3120,RESET,WX3123);
	and 	XG2701 	(WX3118,RESET,WX3121);
	and 	XG2702 	(WX3116,RESET,WX3119);
	and 	XG2703 	(WX3114,RESET,WX3117);
	and 	XG2704 	(WX3112,RESET,WX3115);
	and 	XG2705 	(WX3110,RESET,WX3113);
	and 	XG2706 	(WX3108,RESET,WX3111);
	and 	XG2707 	(WX3106,RESET,WX3109);
	and 	XG2708 	(WX3104,RESET,WX3107);
	and 	XG2709 	(WX3102,RESET,WX3105);
	and 	XG2710 	(WX3100,RESET,WX3103);
	and 	XG2711 	(WX3098,RESET,WX3101);
	and 	XG2712 	(WX3096,RESET,WX3099);
	and 	XG2713 	(WX3094,RESET,WX3097);
	and 	XG2714 	(WX3092,RESET,WX3095);
	and 	XG2715 	(WX3090,RESET,WX3093);
	and 	XG2716 	(WX3088,RESET,WX3091);
	and 	XG2717 	(WX3086,RESET,WX3089);
	and 	XG2718 	(WX3084,RESET,WX3087);
	and 	XG2719 	(WX3082,RESET,WX3085);
	and 	XG2720 	(WX3080,RESET,WX3083);
	and 	XG2721 	(WX3078,RESET,WX3081);
	and 	XG2722 	(WX3076,RESET,WX3079);
	and 	XG2723 	(WX3074,RESET,WX3077);
	and 	XG2724 	(WX3072,RESET,WX3075);
	and 	XG2725 	(WX3070,RESET,WX3073);
	and 	XG2726 	(WX2191,RESET,WX2128);
	and 	XG2727 	(WX2189,RESET,WX2126);
	and 	XG2728 	(WX2187,RESET,WX2124);
	and 	XG2729 	(WX2185,RESET,WX2122);
	and 	XG2730 	(WX2183,RESET,WX2120);
	and 	XG2731 	(WX2181,RESET,WX2118);
	and 	XG2732 	(WX2179,RESET,WX2116);
	and 	XG2733 	(WX2177,RESET,WX2114);
	and 	XG2734 	(WX2175,RESET,WX2112);
	and 	XG2735 	(WX2173,RESET,WX2110);
	and 	XG2736 	(WX2171,RESET,WX2108);
	and 	XG2737 	(WX2169,RESET,WX2106);
	and 	XG2738 	(WX2167,RESET,WX2104);
	and 	XG2739 	(WX2165,RESET,WX2102);
	and 	XG2740 	(WX2163,RESET,WX2100);
	and 	XG2741 	(WX2161,RESET,WX2098);
	and 	XG2742 	(WX2159,RESET,WX2096);
	and 	XG2743 	(WX2157,RESET,WX2094);
	and 	XG2744 	(WX2155,RESET,WX2092);
	and 	XG2745 	(WX2153,RESET,WX2090);
	and 	XG2746 	(WX2151,RESET,WX2088);
	and 	XG2747 	(WX2149,RESET,WX2086);
	and 	XG2748 	(WX2147,RESET,WX2084);
	and 	XG2749 	(WX2145,RESET,WX2082);
	and 	XG2750 	(WX2143,RESET,WX2080);
	and 	XG2751 	(WX2141,RESET,WX2078);
	and 	XG2752 	(WX2139,RESET,WX2076);
	and 	XG2753 	(WX2137,RESET,WX2074);
	and 	XG2754 	(WX2135,RESET,WX2072);
	and 	XG2755 	(WX2133,RESET,WX2070);
	and 	XG2756 	(WX2131,RESET,WX2068);
	and 	XG2757 	(WX2129,RESET,WX2066);
	and 	XG2758 	(WX2127,RESET,WX2064);
	and 	XG2759 	(WX2125,RESET,WX2062);
	and 	XG2760 	(WX2123,RESET,WX2060);
	and 	XG2761 	(WX2121,RESET,WX2058);
	and 	XG2762 	(WX2119,RESET,WX2056);
	and 	XG2763 	(WX2117,RESET,WX2054);
	and 	XG2764 	(WX2115,RESET,WX2052);
	and 	XG2765 	(WX2113,RESET,WX2050);
	and 	XG2766 	(WX2111,RESET,WX2048);
	and 	XG2767 	(WX2109,RESET,WX2046);
	and 	XG2768 	(WX2107,RESET,WX2044);
	and 	XG2769 	(WX2105,RESET,WX2042);
	and 	XG2770 	(WX2103,RESET,WX2040);
	and 	XG2771 	(WX2101,RESET,WX2038);
	and 	XG2772 	(WX2099,RESET,WX2036);
	and 	XG2773 	(WX2097,RESET,WX2034);
	and 	XG2774 	(WX2095,RESET,WX2032);
	and 	XG2775 	(WX2093,RESET,WX2030);
	and 	XG2776 	(WX2091,RESET,WX2028);
	and 	XG2777 	(WX2089,RESET,WX2026);
	and 	XG2778 	(WX2087,RESET,WX2024);
	and 	XG2779 	(WX2085,RESET,WX2022);
	and 	XG2780 	(WX2083,RESET,WX2020);
	and 	XG2781 	(WX2081,RESET,WX2018);
	and 	XG2782 	(WX2079,RESET,WX2016);
	and 	XG2783 	(WX2077,RESET,WX2014);
	and 	XG2784 	(WX2075,RESET,WX2012);
	and 	XG2785 	(WX2073,RESET,WX2010);
	and 	XG2786 	(WX2071,RESET,WX2008);
	and 	XG2787 	(WX2069,RESET,WX2006);
	and 	XG2788 	(WX2067,RESET,WX2004);
	and 	XG2789 	(WX2065,RESET,WX2002);
	and 	XG2790 	(WX2063,RESET,WX2000);
	and 	XG2791 	(WX2061,RESET,WX1998);
	and 	XG2792 	(WX2059,RESET,WX1996);
	and 	XG2793 	(WX2057,RESET,WX1994);
	and 	XG2794 	(WX2055,RESET,WX1992);
	and 	XG2795 	(WX2053,RESET,WX1990);
	and 	XG2796 	(WX2051,RESET,WX1988);
	and 	XG2797 	(WX2049,RESET,WX1986);
	and 	XG2798 	(WX2047,RESET,WX1984);
	and 	XG2799 	(WX2045,RESET,WX1982);
	and 	XG2800 	(WX2043,RESET,WX1980);
	and 	XG2801 	(WX2041,RESET,WX1978);
	and 	XG2802 	(WX2039,RESET,WX1976);
	and 	XG2803 	(WX2037,RESET,WX1974);
	and 	XG2804 	(WX2035,RESET,WX1972);
	and 	XG2805 	(WX2033,RESET,WX1970);
	and 	XG2806 	(WX2031,RESET,WX1968);
	and 	XG2807 	(WX2029,RESET,WX1966);
	and 	XG2808 	(WX2027,RESET,WX1964);
	and 	XG2809 	(WX2025,RESET,WX1962);
	and 	XG2810 	(WX2023,RESET,WX1960);
	and 	XG2811 	(WX2021,RESET,WX1958);
	and 	XG2812 	(WX2019,RESET,WX1956);
	and 	XG2813 	(WX2017,RESET,WX1954);
	and 	XG2814 	(WX2015,RESET,WX1952);
	and 	XG2815 	(WX2013,RESET,WX1950);
	and 	XG2816 	(WX2011,RESET,WX1948);
	and 	XG2817 	(WX2009,RESET,WX1946);
	and 	XG2818 	(WX2007,RESET,WX1944);
	and 	XG2819 	(WX2005,RESET,WX1942);
	and 	XG2820 	(WX2003,RESET,WX1940);
	and 	XG2821 	(WX2001,RESET,WX1938);
	and 	XG2822 	(WX1837,RESET,WX1840);
	and 	XG2823 	(WX1835,RESET,WX1838);
	and 	XG2824 	(WX1833,RESET,WX1836);
	and 	XG2825 	(WX1831,RESET,WX1834);
	and 	XG2826 	(WX1829,RESET,WX1832);
	and 	XG2827 	(WX1827,RESET,WX1830);
	and 	XG2828 	(WX1825,RESET,WX1828);
	and 	XG2829 	(WX1823,RESET,WX1826);
	and 	XG2830 	(WX1821,RESET,WX1824);
	and 	XG2831 	(WX1819,RESET,WX1822);
	and 	XG2832 	(WX1817,RESET,WX1820);
	and 	XG2833 	(WX1815,RESET,WX1818);
	and 	XG2834 	(WX1813,RESET,WX1816);
	and 	XG2835 	(WX1811,RESET,WX1814);
	and 	XG2836 	(WX1809,RESET,WX1812);
	and 	XG2837 	(WX1807,RESET,WX1810);
	and 	XG2838 	(WX1805,RESET,WX1808);
	and 	XG2839 	(WX1803,RESET,WX1806);
	and 	XG2840 	(WX1801,RESET,WX1804);
	and 	XG2841 	(WX1799,RESET,WX1802);
	and 	XG2842 	(WX1797,RESET,WX1800);
	and 	XG2843 	(WX1795,RESET,WX1798);
	and 	XG2844 	(WX1793,RESET,WX1796);
	and 	XG2845 	(WX1791,RESET,WX1794);
	and 	XG2846 	(WX1789,RESET,WX1792);
	and 	XG2847 	(WX1787,RESET,WX1790);
	and 	XG2848 	(WX1785,RESET,WX1788);
	and 	XG2849 	(WX1783,RESET,WX1786);
	and 	XG2850 	(WX1781,RESET,WX1784);
	and 	XG2851 	(WX1779,RESET,WX1782);
	and 	XG2852 	(WX1777,RESET,WX1780);
	and 	XG2853 	(WX898,RESET,WX835);
	and 	XG2854 	(WX896,RESET,WX833);
	and 	XG2855 	(WX894,RESET,WX831);
	and 	XG2856 	(WX892,RESET,WX829);
	and 	XG2857 	(WX890,RESET,WX827);
	and 	XG2858 	(WX888,RESET,WX825);
	and 	XG2859 	(WX886,RESET,WX823);
	and 	XG2860 	(WX884,RESET,WX821);
	and 	XG2861 	(WX882,RESET,WX819);
	and 	XG2862 	(WX880,RESET,WX817);
	and 	XG2863 	(WX878,RESET,WX815);
	and 	XG2864 	(WX876,RESET,WX813);
	and 	XG2865 	(WX874,RESET,WX811);
	and 	XG2866 	(WX872,RESET,WX809);
	and 	XG2867 	(WX870,RESET,WX807);
	and 	XG2868 	(WX868,RESET,WX805);
	and 	XG2869 	(WX866,RESET,WX803);
	and 	XG2870 	(WX864,RESET,WX801);
	and 	XG2871 	(WX862,RESET,WX799);
	and 	XG2872 	(WX860,RESET,WX797);
	and 	XG2873 	(WX858,RESET,WX795);
	and 	XG2874 	(WX856,RESET,WX793);
	and 	XG2875 	(WX854,RESET,WX791);
	and 	XG2876 	(WX852,RESET,WX789);
	and 	XG2877 	(WX850,RESET,WX787);
	and 	XG2878 	(WX848,RESET,WX785);
	and 	XG2879 	(WX846,RESET,WX783);
	and 	XG2880 	(WX844,RESET,WX781);
	and 	XG2881 	(WX842,RESET,WX779);
	and 	XG2882 	(WX840,RESET,WX777);
	and 	XG2883 	(WX838,RESET,WX775);
	and 	XG2884 	(WX836,RESET,WX773);
	and 	XG2885 	(WX834,RESET,WX771);
	and 	XG2886 	(WX832,RESET,WX769);
	and 	XG2887 	(WX830,RESET,WX767);
	and 	XG2888 	(WX828,RESET,WX765);
	and 	XG2889 	(WX826,RESET,WX763);
	and 	XG2890 	(WX824,RESET,WX761);
	and 	XG2891 	(WX822,RESET,WX759);
	and 	XG2892 	(WX820,RESET,WX757);
	and 	XG2893 	(WX818,RESET,WX755);
	and 	XG2894 	(WX816,RESET,WX753);
	and 	XG2895 	(WX814,RESET,WX751);
	and 	XG2896 	(WX812,RESET,WX749);
	and 	XG2897 	(WX810,RESET,WX747);
	and 	XG2898 	(WX808,RESET,WX745);
	and 	XG2899 	(WX806,RESET,WX743);
	and 	XG2900 	(WX804,RESET,WX741);
	and 	XG2901 	(WX802,RESET,WX739);
	and 	XG2902 	(WX800,RESET,WX737);
	and 	XG2903 	(WX798,RESET,WX735);
	and 	XG2904 	(WX796,RESET,WX733);
	and 	XG2905 	(WX794,RESET,WX731);
	and 	XG2906 	(WX792,RESET,WX729);
	and 	XG2907 	(WX790,RESET,WX727);
	and 	XG2908 	(WX788,RESET,WX725);
	and 	XG2909 	(WX786,RESET,WX723);
	and 	XG2910 	(WX784,RESET,WX721);
	and 	XG2911 	(WX782,RESET,WX719);
	and 	XG2912 	(WX780,RESET,WX717);
	and 	XG2913 	(WX778,RESET,WX715);
	and 	XG2914 	(WX776,RESET,WX713);
	and 	XG2915 	(WX774,RESET,WX711);
	and 	XG2916 	(WX772,RESET,WX709);
	and 	XG2917 	(WX770,RESET,WX707);
	and 	XG2918 	(WX768,RESET,WX705);
	and 	XG2919 	(WX766,RESET,WX703);
	and 	XG2920 	(WX764,RESET,WX701);
	and 	XG2921 	(WX762,RESET,WX699);
	and 	XG2922 	(WX760,RESET,WX697);
	and 	XG2923 	(WX758,RESET,WX695);
	and 	XG2924 	(WX756,RESET,WX693);
	and 	XG2925 	(WX754,RESET,WX691);
	and 	XG2926 	(WX752,RESET,WX689);
	and 	XG2927 	(WX750,RESET,WX687);
	and 	XG2928 	(WX748,RESET,WX685);
	and 	XG2929 	(WX746,RESET,WX683);
	and 	XG2930 	(WX744,RESET,WX681);
	and 	XG2931 	(WX742,RESET,WX679);
	and 	XG2932 	(WX740,RESET,WX677);
	and 	XG2933 	(WX738,RESET,WX675);
	and 	XG2934 	(WX736,RESET,WX673);
	and 	XG2935 	(WX734,RESET,WX671);
	and 	XG2936 	(WX732,RESET,WX669);
	and 	XG2937 	(WX730,RESET,WX667);
	and 	XG2938 	(WX728,RESET,WX665);
	and 	XG2939 	(WX726,RESET,WX663);
	and 	XG2940 	(WX724,RESET,WX661);
	and 	XG2941 	(WX722,RESET,WX659);
	and 	XG2942 	(WX720,RESET,WX657);
	and 	XG2943 	(WX718,RESET,WX655);
	and 	XG2944 	(WX716,RESET,WX653);
	and 	XG2945 	(WX714,RESET,WX651);
	and 	XG2946 	(WX712,RESET,WX649);
	and 	XG2947 	(WX710,RESET,WX647);
	and 	XG2948 	(WX708,RESET,WX645);
	and 	XG2949 	(WX544,RESET,WX547);
	and 	XG2950 	(WX542,RESET,WX545);
	and 	XG2951 	(WX540,RESET,WX543);
	and 	XG2952 	(WX538,RESET,WX541);
	and 	XG2953 	(WX536,RESET,WX539);
	and 	XG2954 	(WX534,RESET,WX537);
	and 	XG2955 	(WX532,RESET,WX535);
	and 	XG2956 	(WX530,RESET,WX533);
	and 	XG2957 	(WX528,RESET,WX531);
	and 	XG2958 	(WX526,RESET,WX529);
	and 	XG2959 	(WX524,RESET,WX527);
	and 	XG2960 	(WX522,RESET,WX525);
	and 	XG2961 	(WX520,RESET,WX523);
	and 	XG2962 	(WX518,RESET,WX521);
	and 	XG2963 	(WX516,RESET,WX519);
	and 	XG2964 	(WX514,RESET,WX517);
	and 	XG2965 	(WX512,RESET,WX515);
	and 	XG2966 	(WX510,RESET,WX513);
	and 	XG2967 	(WX508,RESET,WX511);
	and 	XG2968 	(WX506,RESET,WX509);
	and 	XG2969 	(WX504,RESET,WX507);
	and 	XG2970 	(WX502,RESET,WX505);
	and 	XG2971 	(WX500,RESET,WX503);
	and 	XG2972 	(WX498,RESET,WX501);
	and 	XG2973 	(WX496,RESET,WX499);
	and 	XG2974 	(WX494,RESET,WX497);
	and 	XG2975 	(WX492,RESET,WX495);
	and 	XG2976 	(WX490,RESET,WX493);
	and 	XG2977 	(WX488,RESET,WX491);
	and 	XG2978 	(WX486,RESET,WX489);
	and 	XG2979 	(WX484,RESET,WX487);
	not 	XG2980 	(WX483,WX485);
	nand 	XG2981 	(II2003,WX837,WX773);
	nand 	XG2982 	(II2034,WX839,WX775);
	nand 	XG2983 	(II2065,WX841,WX777);
	nand 	XG2984 	(II2096,WX843,WX779);
	nand 	XG2985 	(II2127,WX845,WX781);
	nand 	XG2986 	(II2158,WX847,WX783);
	nand 	XG2987 	(II2189,WX849,WX785);
	nand 	XG2988 	(II2220,WX851,WX787);
	nand 	XG2989 	(II2251,WX853,WX789);
	nand 	XG2990 	(II2282,WX855,WX791);
	nand 	XG2991 	(II2313,WX857,WX793);
	nand 	XG2992 	(II2344,WX859,WX795);
	nand 	XG2993 	(II2375,WX861,WX797);
	nand 	XG2994 	(II2406,WX863,WX799);
	nand 	XG2995 	(II2437,WX865,WX801);
	nand 	XG2996 	(II2468,WX867,WX803);
	nand 	XG2997 	(II2499,WX869,WX805);
	nand 	XG2998 	(II2530,WX871,WX807);
	nand 	XG2999 	(II2561,WX873,WX809);
	nand 	XG3000 	(II2592,WX875,WX811);
	nand 	XG3001 	(II2623,WX877,WX813);
	nand 	XG3002 	(II2654,WX879,WX815);
	nand 	XG3003 	(II2685,WX881,WX817);
	nand 	XG3004 	(II2716,WX883,WX819);
	nand 	XG3005 	(II2747,WX885,WX821);
	nand 	XG3006 	(II2778,WX887,WX823);
	nand 	XG3007 	(II2809,WX889,WX825);
	nand 	XG3008 	(II2840,WX891,WX827);
	nand 	XG3009 	(II2871,WX893,WX829);
	nand 	XG3010 	(II2902,WX895,WX831);
	nand 	XG3011 	(II2933,WX897,WX833);
	nand 	XG3012 	(II2964,WX899,WX835);
	not 	XG3013 	(WX612,WX837);
	not 	XG3014 	(WX613,WX839);
	not 	XG3015 	(WX614,WX841);
	not 	XG3016 	(WX615,WX843);
	not 	XG3017 	(WX616,WX845);
	not 	XG3018 	(WX617,WX847);
	not 	XG3019 	(WX618,WX849);
	not 	XG3020 	(WX619,WX851);
	not 	XG3021 	(WX620,WX853);
	not 	XG3022 	(WX621,WX855);
	not 	XG3023 	(WX622,WX857);
	not 	XG3024 	(WX623,WX859);
	not 	XG3025 	(WX624,WX861);
	not 	XG3026 	(WX625,WX863);
	not 	XG3027 	(WX626,WX865);
	not 	XG3028 	(WX627,WX867);
	not 	XG3029 	(WX628,WX869);
	not 	XG3030 	(WX629,WX871);
	not 	XG3031 	(WX630,WX873);
	not 	XG3032 	(WX631,WX875);
	not 	XG3033 	(WX632,WX877);
	not 	XG3034 	(WX633,WX879);
	not 	XG3035 	(WX634,WX881);
	not 	XG3036 	(WX635,WX883);
	not 	XG3037 	(WX636,WX885);
	not 	XG3038 	(WX637,WX887);
	not 	XG3039 	(WX638,WX889);
	not 	XG3040 	(WX639,WX891);
	not 	XG3041 	(WX640,WX893);
	not 	XG3042 	(WX641,WX895);
	not 	XG3043 	(WX642,WX897);
	not 	XG3044 	(WX643,WX899);
	not 	XG3045 	(WX1776,WX1778);
	nand 	XG3046 	(II6008,WX2130,WX2066);
	nand 	XG3047 	(II6039,WX2132,WX2068);
	nand 	XG3048 	(II6070,WX2134,WX2070);
	nand 	XG3049 	(II6101,WX2136,WX2072);
	nand 	XG3050 	(II6132,WX2138,WX2074);
	nand 	XG3051 	(II6163,WX2140,WX2076);
	nand 	XG3052 	(II6194,WX2142,WX2078);
	nand 	XG3053 	(II6225,WX2144,WX2080);
	nand 	XG3054 	(II6256,WX2146,WX2082);
	nand 	XG3055 	(II6287,WX2148,WX2084);
	nand 	XG3056 	(II6318,WX2150,WX2086);
	nand 	XG3057 	(II6349,WX2152,WX2088);
	nand 	XG3058 	(II6380,WX2154,WX2090);
	nand 	XG3059 	(II6411,WX2156,WX2092);
	nand 	XG3060 	(II6442,WX2158,WX2094);
	nand 	XG3061 	(II6473,WX2160,WX2096);
	nand 	XG3062 	(II6504,WX2162,WX2098);
	nand 	XG3063 	(II6535,WX2164,WX2100);
	nand 	XG3064 	(II6566,WX2166,WX2102);
	nand 	XG3065 	(II6597,WX2168,WX2104);
	nand 	XG3066 	(II6628,WX2170,WX2106);
	nand 	XG3067 	(II6659,WX2172,WX2108);
	nand 	XG3068 	(II6690,WX2174,WX2110);
	nand 	XG3069 	(II6721,WX2176,WX2112);
	nand 	XG3070 	(II6752,WX2178,WX2114);
	nand 	XG3071 	(II6783,WX2180,WX2116);
	nand 	XG3072 	(II6814,WX2182,WX2118);
	nand 	XG3073 	(II6845,WX2184,WX2120);
	nand 	XG3074 	(II6876,WX2186,WX2122);
	nand 	XG3075 	(II6907,WX2188,WX2124);
	nand 	XG3076 	(II6938,WX2190,WX2126);
	nand 	XG3077 	(II6969,WX2192,WX2128);
	not 	XG3078 	(WX1905,WX2130);
	not 	XG3079 	(WX1906,WX2132);
	not 	XG3080 	(WX1907,WX2134);
	not 	XG3081 	(WX1908,WX2136);
	not 	XG3082 	(WX1909,WX2138);
	not 	XG3083 	(WX1910,WX2140);
	not 	XG3084 	(WX1911,WX2142);
	not 	XG3085 	(WX1912,WX2144);
	not 	XG3086 	(WX1913,WX2146);
	not 	XG3087 	(WX1914,WX2148);
	not 	XG3088 	(WX1915,WX2150);
	not 	XG3089 	(WX1916,WX2152);
	not 	XG3090 	(WX1917,WX2154);
	not 	XG3091 	(WX1918,WX2156);
	not 	XG3092 	(WX1919,WX2158);
	not 	XG3093 	(WX1920,WX2160);
	not 	XG3094 	(WX1921,WX2162);
	not 	XG3095 	(WX1922,WX2164);
	not 	XG3096 	(WX1923,WX2166);
	not 	XG3097 	(WX1924,WX2168);
	not 	XG3098 	(WX1925,WX2170);
	not 	XG3099 	(WX1926,WX2172);
	not 	XG3100 	(WX1927,WX2174);
	not 	XG3101 	(WX1928,WX2176);
	not 	XG3102 	(WX1929,WX2178);
	not 	XG3103 	(WX1930,WX2180);
	not 	XG3104 	(WX1931,WX2182);
	not 	XG3105 	(WX1932,WX2184);
	not 	XG3106 	(WX1933,WX2186);
	not 	XG3107 	(WX1934,WX2188);
	not 	XG3108 	(WX1935,WX2190);
	not 	XG3109 	(WX1936,WX2192);
	not 	XG3110 	(WX3069,WX3071);
	nand 	XG3111 	(II10013,WX3423,WX3359);
	nand 	XG3112 	(II10044,WX3425,WX3361);
	nand 	XG3113 	(II10075,WX3427,WX3363);
	nand 	XG3114 	(II10106,WX3429,WX3365);
	nand 	XG3115 	(II10137,WX3431,WX3367);
	nand 	XG3116 	(II10168,WX3433,WX3369);
	nand 	XG3117 	(II10199,WX3435,WX3371);
	nand 	XG3118 	(II10230,WX3437,WX3373);
	nand 	XG3119 	(II10261,WX3439,WX3375);
	nand 	XG3120 	(II10292,WX3441,WX3377);
	nand 	XG3121 	(II10323,WX3443,WX3379);
	nand 	XG3122 	(II10354,WX3445,WX3381);
	nand 	XG3123 	(II10385,WX3447,WX3383);
	nand 	XG3124 	(II10416,WX3449,WX3385);
	nand 	XG3125 	(II10447,WX3451,WX3387);
	nand 	XG3126 	(II10478,WX3453,WX3389);
	nand 	XG3127 	(II10509,WX3455,WX3391);
	nand 	XG3128 	(II10540,WX3457,WX3393);
	nand 	XG3129 	(II10571,WX3459,WX3395);
	nand 	XG3130 	(II10602,WX3461,WX3397);
	nand 	XG3131 	(II10633,WX3463,WX3399);
	nand 	XG3132 	(II10664,WX3465,WX3401);
	nand 	XG3133 	(II10695,WX3467,WX3403);
	nand 	XG3134 	(II10726,WX3469,WX3405);
	nand 	XG3135 	(II10757,WX3471,WX3407);
	nand 	XG3136 	(II10788,WX3473,WX3409);
	nand 	XG3137 	(II10819,WX3475,WX3411);
	nand 	XG3138 	(II10850,WX3477,WX3413);
	nand 	XG3139 	(II10881,WX3479,WX3415);
	nand 	XG3140 	(II10912,WX3481,WX3417);
	nand 	XG3141 	(II10943,WX3483,WX3419);
	nand 	XG3142 	(II10974,WX3485,WX3421);
	not 	XG3143 	(WX3198,WX3423);
	not 	XG3144 	(WX3199,WX3425);
	not 	XG3145 	(WX3200,WX3427);
	not 	XG3146 	(WX3201,WX3429);
	not 	XG3147 	(WX3202,WX3431);
	not 	XG3148 	(WX3203,WX3433);
	not 	XG3149 	(WX3204,WX3435);
	not 	XG3150 	(WX3205,WX3437);
	not 	XG3151 	(WX3206,WX3439);
	not 	XG3152 	(WX3207,WX3441);
	not 	XG3153 	(WX3208,WX3443);
	not 	XG3154 	(WX3209,WX3445);
	not 	XG3155 	(WX3210,WX3447);
	not 	XG3156 	(WX3211,WX3449);
	not 	XG3157 	(WX3212,WX3451);
	not 	XG3158 	(WX3213,WX3453);
	not 	XG3159 	(WX3214,WX3455);
	not 	XG3160 	(WX3215,WX3457);
	not 	XG3161 	(WX3216,WX3459);
	not 	XG3162 	(WX3217,WX3461);
	not 	XG3163 	(WX3218,WX3463);
	not 	XG3164 	(WX3219,WX3465);
	not 	XG3165 	(WX3220,WX3467);
	not 	XG3166 	(WX3221,WX3469);
	not 	XG3167 	(WX3222,WX3471);
	not 	XG3168 	(WX3223,WX3473);
	not 	XG3169 	(WX3224,WX3475);
	not 	XG3170 	(WX3225,WX3477);
	not 	XG3171 	(WX3226,WX3479);
	not 	XG3172 	(WX3227,WX3481);
	not 	XG3173 	(WX3228,WX3483);
	not 	XG3174 	(WX3229,WX3485);
	not 	XG3175 	(WX4362,WX4364);
	nand 	XG3176 	(II14018,WX4716,WX4652);
	nand 	XG3177 	(II14049,WX4718,WX4654);
	nand 	XG3178 	(II14080,WX4720,WX4656);
	nand 	XG3179 	(II14111,WX4722,WX4658);
	nand 	XG3180 	(II14142,WX4724,WX4660);
	nand 	XG3181 	(II14173,WX4726,WX4662);
	nand 	XG3182 	(II14204,WX4728,WX4664);
	nand 	XG3183 	(II14235,WX4730,WX4666);
	nand 	XG3184 	(II14266,WX4732,WX4668);
	nand 	XG3185 	(II14297,WX4734,WX4670);
	nand 	XG3186 	(II14328,WX4736,WX4672);
	nand 	XG3187 	(II14359,WX4738,WX4674);
	nand 	XG3188 	(II14390,WX4740,WX4676);
	nand 	XG3189 	(II14421,WX4742,WX4678);
	nand 	XG3190 	(II14452,WX4744,WX4680);
	nand 	XG3191 	(II14483,WX4746,WX4682);
	nand 	XG3192 	(II14514,WX4748,WX4684);
	nand 	XG3193 	(II14545,WX4750,WX4686);
	nand 	XG3194 	(II14576,WX4752,WX4688);
	nand 	XG3195 	(II14607,WX4754,WX4690);
	nand 	XG3196 	(II14638,WX4756,WX4692);
	nand 	XG3197 	(II14669,WX4758,WX4694);
	nand 	XG3198 	(II14700,WX4760,WX4696);
	nand 	XG3199 	(II14731,WX4762,WX4698);
	nand 	XG3200 	(II14762,WX4764,WX4700);
	nand 	XG3201 	(II14793,WX4766,WX4702);
	nand 	XG3202 	(II14824,WX4768,WX4704);
	nand 	XG3203 	(II14855,WX4770,WX4706);
	nand 	XG3204 	(II14886,WX4772,WX4708);
	nand 	XG3205 	(II14917,WX4774,WX4710);
	nand 	XG3206 	(II14948,WX4776,WX4712);
	nand 	XG3207 	(II14979,WX4778,WX4714);
	not 	XG3208 	(WX4491,WX4716);
	not 	XG3209 	(WX4492,WX4718);
	not 	XG3210 	(WX4493,WX4720);
	not 	XG3211 	(WX4494,WX4722);
	not 	XG3212 	(WX4495,WX4724);
	not 	XG3213 	(WX4496,WX4726);
	not 	XG3214 	(WX4497,WX4728);
	not 	XG3215 	(WX4498,WX4730);
	not 	XG3216 	(WX4499,WX4732);
	not 	XG3217 	(WX4500,WX4734);
	not 	XG3218 	(WX4501,WX4736);
	not 	XG3219 	(WX4502,WX4738);
	not 	XG3220 	(WX4503,WX4740);
	not 	XG3221 	(WX4504,WX4742);
	not 	XG3222 	(WX4505,WX4744);
	not 	XG3223 	(WX4506,WX4746);
	not 	XG3224 	(WX4507,WX4748);
	not 	XG3225 	(WX4508,WX4750);
	not 	XG3226 	(WX4509,WX4752);
	not 	XG3227 	(WX4510,WX4754);
	not 	XG3228 	(WX4511,WX4756);
	not 	XG3229 	(WX4512,WX4758);
	not 	XG3230 	(WX4513,WX4760);
	not 	XG3231 	(WX4514,WX4762);
	not 	XG3232 	(WX4515,WX4764);
	not 	XG3233 	(WX4516,WX4766);
	not 	XG3234 	(WX4517,WX4768);
	not 	XG3235 	(WX4518,WX4770);
	not 	XG3236 	(WX4519,WX4772);
	not 	XG3237 	(WX4520,WX4774);
	not 	XG3238 	(WX4521,WX4776);
	not 	XG3239 	(WX4522,WX4778);
	not 	XG3240 	(WX5655,WX5657);
	nand 	XG3241 	(II18023,WX6009,WX5945);
	nand 	XG3242 	(II18054,WX6011,WX5947);
	nand 	XG3243 	(II18085,WX6013,WX5949);
	nand 	XG3244 	(II18116,WX6015,WX5951);
	nand 	XG3245 	(II18147,WX6017,WX5953);
	nand 	XG3246 	(II18178,WX6019,WX5955);
	nand 	XG3247 	(II18209,WX6021,WX5957);
	nand 	XG3248 	(II18240,WX6023,WX5959);
	nand 	XG3249 	(II18271,WX6025,WX5961);
	nand 	XG3250 	(II18302,WX6027,WX5963);
	nand 	XG3251 	(II18333,WX6029,WX5965);
	nand 	XG3252 	(II18364,WX6031,WX5967);
	nand 	XG3253 	(II18395,WX6033,WX5969);
	nand 	XG3254 	(II18426,WX6035,WX5971);
	nand 	XG3255 	(II18457,WX6037,WX5973);
	nand 	XG3256 	(II18488,WX6039,WX5975);
	nand 	XG3257 	(II18519,WX6041,WX5977);
	nand 	XG3258 	(II18550,WX6043,WX5979);
	nand 	XG3259 	(II18581,WX6045,WX5981);
	nand 	XG3260 	(II18612,WX6047,WX5983);
	nand 	XG3261 	(II18643,WX6049,WX5985);
	nand 	XG3262 	(II18674,WX6051,WX5987);
	nand 	XG3263 	(II18705,WX6053,WX5989);
	nand 	XG3264 	(II18736,WX6055,WX5991);
	nand 	XG3265 	(II18767,WX6057,WX5993);
	nand 	XG3266 	(II18798,WX6059,WX5995);
	nand 	XG3267 	(II18829,WX6061,WX5997);
	nand 	XG3268 	(II18860,WX6063,WX5999);
	nand 	XG3269 	(II18891,WX6065,WX6001);
	nand 	XG3270 	(II18922,WX6067,WX6003);
	nand 	XG3271 	(II18953,WX6069,WX6005);
	nand 	XG3272 	(II18984,WX6071,WX6007);
	not 	XG3273 	(WX5784,WX6009);
	not 	XG3274 	(WX5785,WX6011);
	not 	XG3275 	(WX5786,WX6013);
	not 	XG3276 	(WX5787,WX6015);
	not 	XG3277 	(WX5788,WX6017);
	not 	XG3278 	(WX5789,WX6019);
	not 	XG3279 	(WX5790,WX6021);
	not 	XG3280 	(WX5791,WX6023);
	not 	XG3281 	(WX5792,WX6025);
	not 	XG3282 	(WX5793,WX6027);
	not 	XG3283 	(WX5794,WX6029);
	not 	XG3284 	(WX5795,WX6031);
	not 	XG3285 	(WX5796,WX6033);
	not 	XG3286 	(WX5797,WX6035);
	not 	XG3287 	(WX5798,WX6037);
	not 	XG3288 	(WX5799,WX6039);
	not 	XG3289 	(WX5800,WX6041);
	not 	XG3290 	(WX5801,WX6043);
	not 	XG3291 	(WX5802,WX6045);
	not 	XG3292 	(WX5803,WX6047);
	not 	XG3293 	(WX5804,WX6049);
	not 	XG3294 	(WX5805,WX6051);
	not 	XG3295 	(WX5806,WX6053);
	not 	XG3296 	(WX5807,WX6055);
	not 	XG3297 	(WX5808,WX6057);
	not 	XG3298 	(WX5809,WX6059);
	not 	XG3299 	(WX5810,WX6061);
	not 	XG3300 	(WX5811,WX6063);
	not 	XG3301 	(WX5812,WX6065);
	not 	XG3302 	(WX5813,WX6067);
	not 	XG3303 	(WX5814,WX6069);
	not 	XG3304 	(WX5815,WX6071);
	not 	XG3305 	(WX6948,WX6950);
	nand 	XG3306 	(II22028,WX7302,WX7238);
	nand 	XG3307 	(II22059,WX7304,WX7240);
	nand 	XG3308 	(II22090,WX7306,WX7242);
	nand 	XG3309 	(II22121,WX7308,WX7244);
	nand 	XG3310 	(II22152,WX7310,WX7246);
	nand 	XG3311 	(II22183,WX7312,WX7248);
	nand 	XG3312 	(II22214,WX7314,WX7250);
	nand 	XG3313 	(II22245,WX7316,WX7252);
	nand 	XG3314 	(II22276,WX7318,WX7254);
	nand 	XG3315 	(II22307,WX7320,WX7256);
	nand 	XG3316 	(II22338,WX7322,WX7258);
	nand 	XG3317 	(II22369,WX7324,WX7260);
	nand 	XG3318 	(II22400,WX7326,WX7262);
	nand 	XG3319 	(II22431,WX7328,WX7264);
	nand 	XG3320 	(II22462,WX7330,WX7266);
	nand 	XG3321 	(II22493,WX7332,WX7268);
	nand 	XG3322 	(II22524,WX7334,WX7270);
	nand 	XG3323 	(II22555,WX7336,WX7272);
	nand 	XG3324 	(II22586,WX7338,WX7274);
	nand 	XG3325 	(II22617,WX7340,WX7276);
	nand 	XG3326 	(II22648,WX7342,WX7278);
	nand 	XG3327 	(II22679,WX7344,WX7280);
	nand 	XG3328 	(II22710,WX7346,WX7282);
	nand 	XG3329 	(II22741,WX7348,WX7284);
	nand 	XG3330 	(II22772,WX7350,WX7286);
	nand 	XG3331 	(II22803,WX7352,WX7288);
	nand 	XG3332 	(II22834,WX7354,WX7290);
	nand 	XG3333 	(II22865,WX7356,WX7292);
	nand 	XG3334 	(II22896,WX7358,WX7294);
	nand 	XG3335 	(II22927,WX7360,WX7296);
	nand 	XG3336 	(II22958,WX7362,WX7298);
	nand 	XG3337 	(II22989,WX7364,WX7300);
	not 	XG3338 	(WX7077,WX7302);
	not 	XG3339 	(WX7078,WX7304);
	not 	XG3340 	(WX7079,WX7306);
	not 	XG3341 	(WX7080,WX7308);
	not 	XG3342 	(WX7081,WX7310);
	not 	XG3343 	(WX7082,WX7312);
	not 	XG3344 	(WX7083,WX7314);
	not 	XG3345 	(WX7084,WX7316);
	not 	XG3346 	(WX7085,WX7318);
	not 	XG3347 	(WX7086,WX7320);
	not 	XG3348 	(WX7087,WX7322);
	not 	XG3349 	(WX7088,WX7324);
	not 	XG3350 	(WX7089,WX7326);
	not 	XG3351 	(WX7090,WX7328);
	not 	XG3352 	(WX7091,WX7330);
	not 	XG3353 	(WX7092,WX7332);
	not 	XG3354 	(WX7093,WX7334);
	not 	XG3355 	(WX7094,WX7336);
	not 	XG3356 	(WX7095,WX7338);
	not 	XG3357 	(WX7096,WX7340);
	not 	XG3358 	(WX7097,WX7342);
	not 	XG3359 	(WX7098,WX7344);
	not 	XG3360 	(WX7099,WX7346);
	not 	XG3361 	(WX7100,WX7348);
	not 	XG3362 	(WX7101,WX7350);
	not 	XG3363 	(WX7102,WX7352);
	not 	XG3364 	(WX7103,WX7354);
	not 	XG3365 	(WX7104,WX7356);
	not 	XG3366 	(WX7105,WX7358);
	not 	XG3367 	(WX7106,WX7360);
	not 	XG3368 	(WX7107,WX7362);
	not 	XG3369 	(WX7108,WX7364);
	not 	XG3370 	(WX8241,WX8243);
	nand 	XG3371 	(II26033,WX8595,WX8531);
	nand 	XG3372 	(II26064,WX8597,WX8533);
	nand 	XG3373 	(II26095,WX8599,WX8535);
	nand 	XG3374 	(II26126,WX8601,WX8537);
	nand 	XG3375 	(II26157,WX8603,WX8539);
	nand 	XG3376 	(II26188,WX8605,WX8541);
	nand 	XG3377 	(II26219,WX8607,WX8543);
	nand 	XG3378 	(II26250,WX8609,WX8545);
	nand 	XG3379 	(II26281,WX8611,WX8547);
	nand 	XG3380 	(II26312,WX8613,WX8549);
	nand 	XG3381 	(II26343,WX8615,WX8551);
	nand 	XG3382 	(II26374,WX8617,WX8553);
	nand 	XG3383 	(II26405,WX8619,WX8555);
	nand 	XG3384 	(II26436,WX8621,WX8557);
	nand 	XG3385 	(II26467,WX8623,WX8559);
	nand 	XG3386 	(II26498,WX8625,WX8561);
	nand 	XG3387 	(II26529,WX8627,WX8563);
	nand 	XG3388 	(II26560,WX8629,WX8565);
	nand 	XG3389 	(II26591,WX8631,WX8567);
	nand 	XG3390 	(II26622,WX8633,WX8569);
	nand 	XG3391 	(II26653,WX8635,WX8571);
	nand 	XG3392 	(II26684,WX8637,WX8573);
	nand 	XG3393 	(II26715,WX8639,WX8575);
	nand 	XG3394 	(II26746,WX8641,WX8577);
	nand 	XG3395 	(II26777,WX8643,WX8579);
	nand 	XG3396 	(II26808,WX8645,WX8581);
	nand 	XG3397 	(II26839,WX8647,WX8583);
	nand 	XG3398 	(II26870,WX8649,WX8585);
	nand 	XG3399 	(II26901,WX8651,WX8587);
	nand 	XG3400 	(II26932,WX8653,WX8589);
	nand 	XG3401 	(II26963,WX8655,WX8591);
	nand 	XG3402 	(II26994,WX8657,WX8593);
	not 	XG3403 	(WX8370,WX8595);
	not 	XG3404 	(WX8371,WX8597);
	not 	XG3405 	(WX8372,WX8599);
	not 	XG3406 	(WX8373,WX8601);
	not 	XG3407 	(WX8374,WX8603);
	not 	XG3408 	(WX8375,WX8605);
	not 	XG3409 	(WX8376,WX8607);
	not 	XG3410 	(WX8377,WX8609);
	not 	XG3411 	(WX8378,WX8611);
	not 	XG3412 	(WX8379,WX8613);
	not 	XG3413 	(WX8380,WX8615);
	not 	XG3414 	(WX8381,WX8617);
	not 	XG3415 	(WX8382,WX8619);
	not 	XG3416 	(WX8383,WX8621);
	not 	XG3417 	(WX8384,WX8623);
	not 	XG3418 	(WX8385,WX8625);
	not 	XG3419 	(WX8386,WX8627);
	not 	XG3420 	(WX8387,WX8629);
	not 	XG3421 	(WX8388,WX8631);
	not 	XG3422 	(WX8389,WX8633);
	not 	XG3423 	(WX8390,WX8635);
	not 	XG3424 	(WX8391,WX8637);
	not 	XG3425 	(WX8392,WX8639);
	not 	XG3426 	(WX8393,WX8641);
	not 	XG3427 	(WX8394,WX8643);
	not 	XG3428 	(WX8395,WX8645);
	not 	XG3429 	(WX8396,WX8647);
	not 	XG3430 	(WX8397,WX8649);
	not 	XG3431 	(WX8398,WX8651);
	not 	XG3432 	(WX8399,WX8653);
	not 	XG3433 	(WX8400,WX8655);
	not 	XG3434 	(WX8401,WX8657);
	not 	XG3435 	(WX9534,WX9536);
	nand 	XG3436 	(II30038,WX9888,WX9824);
	nand 	XG3437 	(II30069,WX9890,WX9826);
	nand 	XG3438 	(II30100,WX9892,WX9828);
	nand 	XG3439 	(II30131,WX9894,WX9830);
	nand 	XG3440 	(II30162,WX9896,WX9832);
	nand 	XG3441 	(II30193,WX9898,WX9834);
	nand 	XG3442 	(II30224,WX9900,WX9836);
	nand 	XG3443 	(II30255,WX9902,WX9838);
	nand 	XG3444 	(II30286,WX9904,WX9840);
	nand 	XG3445 	(II30317,WX9906,WX9842);
	nand 	XG3446 	(II30348,WX9908,WX9844);
	nand 	XG3447 	(II30379,WX9910,WX9846);
	nand 	XG3448 	(II30410,WX9912,WX9848);
	nand 	XG3449 	(II30441,WX9914,WX9850);
	nand 	XG3450 	(II30472,WX9916,WX9852);
	nand 	XG3451 	(II30503,WX9918,WX9854);
	nand 	XG3452 	(II30534,WX9920,WX9856);
	nand 	XG3453 	(II30565,WX9922,WX9858);
	nand 	XG3454 	(II30596,WX9924,WX9860);
	nand 	XG3455 	(II30627,WX9926,WX9862);
	nand 	XG3456 	(II30658,WX9928,WX9864);
	nand 	XG3457 	(II30689,WX9930,WX9866);
	nand 	XG3458 	(II30720,WX9932,WX9868);
	nand 	XG3459 	(II30751,WX9934,WX9870);
	nand 	XG3460 	(II30782,WX9936,WX9872);
	nand 	XG3461 	(II30813,WX9938,WX9874);
	nand 	XG3462 	(II30844,WX9940,WX9876);
	nand 	XG3463 	(II30875,WX9942,WX9878);
	nand 	XG3464 	(II30906,WX9944,WX9880);
	nand 	XG3465 	(II30937,WX9946,WX9882);
	nand 	XG3466 	(II30968,WX9948,WX9884);
	nand 	XG3467 	(II30999,WX9950,WX9886);
	not 	XG3468 	(WX9663,WX9888);
	not 	XG3469 	(WX9664,WX9890);
	not 	XG3470 	(WX9665,WX9892);
	not 	XG3471 	(WX9666,WX9894);
	not 	XG3472 	(WX9667,WX9896);
	not 	XG3473 	(WX9668,WX9898);
	not 	XG3474 	(WX9669,WX9900);
	not 	XG3475 	(WX9670,WX9902);
	not 	XG3476 	(WX9671,WX9904);
	not 	XG3477 	(WX9672,WX9906);
	not 	XG3478 	(WX9673,WX9908);
	not 	XG3479 	(WX9674,WX9910);
	not 	XG3480 	(WX9675,WX9912);
	not 	XG3481 	(WX9676,WX9914);
	not 	XG3482 	(WX9677,WX9916);
	not 	XG3483 	(WX9678,WX9918);
	not 	XG3484 	(WX9679,WX9920);
	not 	XG3485 	(WX9680,WX9922);
	not 	XG3486 	(WX9681,WX9924);
	not 	XG3487 	(WX9682,WX9926);
	not 	XG3488 	(WX9683,WX9928);
	not 	XG3489 	(WX9684,WX9930);
	not 	XG3490 	(WX9685,WX9932);
	not 	XG3491 	(WX9686,WX9934);
	not 	XG3492 	(WX9687,WX9936);
	not 	XG3493 	(WX9688,WX9938);
	not 	XG3494 	(WX9689,WX9940);
	not 	XG3495 	(WX9690,WX9942);
	not 	XG3496 	(WX9691,WX9944);
	not 	XG3497 	(WX9692,WX9946);
	not 	XG3498 	(WX9693,WX9948);
	not 	XG3499 	(WX9694,WX9950);
	not 	XG3500 	(WX10827,WX10829);
	nand 	XG3501 	(II34043,WX11181,WX11117);
	nand 	XG3502 	(II34074,WX11183,WX11119);
	nand 	XG3503 	(II34105,WX11185,WX11121);
	nand 	XG3504 	(II34136,WX11187,WX11123);
	nand 	XG3505 	(II34167,WX11189,WX11125);
	nand 	XG3506 	(II34198,WX11191,WX11127);
	nand 	XG3507 	(II34229,WX11193,WX11129);
	nand 	XG3508 	(II34260,WX11195,WX11131);
	nand 	XG3509 	(II34291,WX11197,WX11133);
	nand 	XG3510 	(II34322,WX11199,WX11135);
	nand 	XG3511 	(II34353,WX11201,WX11137);
	nand 	XG3512 	(II34384,WX11203,WX11139);
	nand 	XG3513 	(II34415,WX11205,WX11141);
	nand 	XG3514 	(II34446,WX11207,WX11143);
	nand 	XG3515 	(II34477,WX11209,WX11145);
	nand 	XG3516 	(II34508,WX11211,WX11147);
	nand 	XG3517 	(II34539,WX11213,WX11149);
	nand 	XG3518 	(II34570,WX11215,WX11151);
	nand 	XG3519 	(II34601,WX11217,WX11153);
	nand 	XG3520 	(II34632,WX11219,WX11155);
	nand 	XG3521 	(II34663,WX11221,WX11157);
	nand 	XG3522 	(II34694,WX11223,WX11159);
	nand 	XG3523 	(II34725,WX11225,WX11161);
	nand 	XG3524 	(II34756,WX11227,WX11163);
	nand 	XG3525 	(II34787,WX11229,WX11165);
	nand 	XG3526 	(II34818,WX11231,WX11167);
	nand 	XG3527 	(II34849,WX11233,WX11169);
	nand 	XG3528 	(II34880,WX11235,WX11171);
	nand 	XG3529 	(II34911,WX11237,WX11173);
	nand 	XG3530 	(II34942,WX11239,WX11175);
	nand 	XG3531 	(II34973,WX11241,WX11177);
	nand 	XG3532 	(II35004,WX11243,WX11179);
	not 	XG3533 	(WX10956,WX11181);
	not 	XG3534 	(WX10957,WX11183);
	not 	XG3535 	(WX10958,WX11185);
	not 	XG3536 	(WX10959,WX11187);
	not 	XG3537 	(WX10960,WX11189);
	not 	XG3538 	(WX10961,WX11191);
	not 	XG3539 	(WX10962,WX11193);
	not 	XG3540 	(WX10963,WX11195);
	not 	XG3541 	(WX10964,WX11197);
	not 	XG3542 	(WX10965,WX11199);
	not 	XG3543 	(WX10966,WX11201);
	not 	XG3544 	(WX10967,WX11203);
	not 	XG3545 	(WX10968,WX11205);
	not 	XG3546 	(WX10969,WX11207);
	not 	XG3547 	(WX10970,WX11209);
	not 	XG3548 	(WX10971,WX11211);
	not 	XG3549 	(WX10972,WX11213);
	not 	XG3550 	(WX10973,WX11215);
	not 	XG3551 	(WX10974,WX11217);
	not 	XG3552 	(WX10975,WX11219);
	not 	XG3553 	(WX10976,WX11221);
	not 	XG3554 	(WX10977,WX11223);
	not 	XG3555 	(WX10978,WX11225);
	not 	XG3556 	(WX10979,WX11227);
	not 	XG3557 	(WX10980,WX11229);
	not 	XG3558 	(WX10981,WX11231);
	not 	XG3559 	(WX10982,WX11233);
	not 	XG3560 	(WX10983,WX11235);
	not 	XG3561 	(WX10984,WX11237);
	not 	XG3562 	(WX10985,WX11239);
	not 	XG3563 	(WX10986,WX11241);
	not 	XG3564 	(WX10987,WX11243);
	not 	XG3565 	(WX10815,WX11347);
	not 	XG3566 	(WX10801,WX11347);
	not 	XG3567 	(WX10787,WX11347);
	not 	XG3568 	(WX10773,WX11347);
	not 	XG3569 	(WX10759,WX11347);
	not 	XG3570 	(WX10745,WX11347);
	not 	XG3571 	(WX10731,WX11347);
	not 	XG3572 	(WX10717,WX11347);
	not 	XG3573 	(WX10703,WX11347);
	not 	XG3574 	(WX10689,WX11347);
	not 	XG3575 	(WX10675,WX11347);
	not 	XG3576 	(WX10661,WX11347);
	not 	XG3577 	(WX10647,WX11347);
	not 	XG3578 	(WX10633,WX11347);
	not 	XG3579 	(WX10619,WX11347);
	not 	XG3580 	(WX10605,WX11347);
	not 	XG3581 	(WX10591,WX11347);
	not 	XG3582 	(WX10577,WX11347);
	not 	XG3583 	(WX10563,WX11347);
	not 	XG3584 	(WX10549,WX11347);
	not 	XG3585 	(WX10535,WX11347);
	not 	XG3586 	(WX10521,WX11347);
	not 	XG3587 	(WX10507,WX11347);
	not 	XG3588 	(WX10493,WX11347);
	not 	XG3589 	(WX10479,WX11347);
	not 	XG3590 	(WX10465,WX11347);
	not 	XG3591 	(WX10451,WX11347);
	not 	XG3592 	(WX10437,WX11347);
	not 	XG3593 	(WX10423,WX11347);
	not 	XG3594 	(WX10409,WX11347);
	not 	XG3595 	(WX10395,WX11347);
	not 	XG3596 	(WX10381,WX11347);
	not 	XG3597 	(WX9522,WX10054);
	not 	XG3598 	(WX9508,WX10054);
	not 	XG3599 	(WX9494,WX10054);
	not 	XG3600 	(WX9480,WX10054);
	not 	XG3601 	(WX9466,WX10054);
	not 	XG3602 	(WX9452,WX10054);
	not 	XG3603 	(WX9438,WX10054);
	not 	XG3604 	(WX9424,WX10054);
	not 	XG3605 	(WX9410,WX10054);
	not 	XG3606 	(WX9396,WX10054);
	not 	XG3607 	(WX9382,WX10054);
	not 	XG3608 	(WX9368,WX10054);
	not 	XG3609 	(WX9354,WX10054);
	not 	XG3610 	(WX9340,WX10054);
	not 	XG3611 	(WX9326,WX10054);
	not 	XG3612 	(WX9312,WX10054);
	not 	XG3613 	(WX9298,WX10054);
	not 	XG3614 	(WX9284,WX10054);
	not 	XG3615 	(WX9270,WX10054);
	not 	XG3616 	(WX9256,WX10054);
	not 	XG3617 	(WX9242,WX10054);
	not 	XG3618 	(WX9228,WX10054);
	not 	XG3619 	(WX9214,WX10054);
	not 	XG3620 	(WX9200,WX10054);
	not 	XG3621 	(WX9186,WX10054);
	not 	XG3622 	(WX9172,WX10054);
	not 	XG3623 	(WX9158,WX10054);
	not 	XG3624 	(WX9144,WX10054);
	not 	XG3625 	(WX9130,WX10054);
	not 	XG3626 	(WX9116,WX10054);
	not 	XG3627 	(WX9102,WX10054);
	not 	XG3628 	(WX9088,WX10054);
	not 	XG3629 	(WX8229,WX8761);
	not 	XG3630 	(WX8215,WX8761);
	not 	XG3631 	(WX8201,WX8761);
	not 	XG3632 	(WX8187,WX8761);
	not 	XG3633 	(WX8173,WX8761);
	not 	XG3634 	(WX8159,WX8761);
	not 	XG3635 	(WX8145,WX8761);
	not 	XG3636 	(WX8131,WX8761);
	not 	XG3637 	(WX8117,WX8761);
	not 	XG3638 	(WX8103,WX8761);
	not 	XG3639 	(WX8089,WX8761);
	not 	XG3640 	(WX8075,WX8761);
	not 	XG3641 	(WX8061,WX8761);
	not 	XG3642 	(WX8047,WX8761);
	not 	XG3643 	(WX8033,WX8761);
	not 	XG3644 	(WX8019,WX8761);
	not 	XG3645 	(WX8005,WX8761);
	not 	XG3646 	(WX7991,WX8761);
	not 	XG3647 	(WX7977,WX8761);
	not 	XG3648 	(WX7963,WX8761);
	not 	XG3649 	(WX7949,WX8761);
	not 	XG3650 	(WX7935,WX8761);
	not 	XG3651 	(WX7921,WX8761);
	not 	XG3652 	(WX7907,WX8761);
	not 	XG3653 	(WX7893,WX8761);
	not 	XG3654 	(WX7879,WX8761);
	not 	XG3655 	(WX7865,WX8761);
	not 	XG3656 	(WX7851,WX8761);
	not 	XG3657 	(WX7837,WX8761);
	not 	XG3658 	(WX7823,WX8761);
	not 	XG3659 	(WX7809,WX8761);
	not 	XG3660 	(WX7795,WX8761);
	not 	XG3661 	(WX6936,WX7468);
	not 	XG3662 	(WX6922,WX7468);
	not 	XG3663 	(WX6908,WX7468);
	not 	XG3664 	(WX6894,WX7468);
	not 	XG3665 	(WX6880,WX7468);
	not 	XG3666 	(WX6866,WX7468);
	not 	XG3667 	(WX6852,WX7468);
	not 	XG3668 	(WX6838,WX7468);
	not 	XG3669 	(WX6824,WX7468);
	not 	XG3670 	(WX6810,WX7468);
	not 	XG3671 	(WX6796,WX7468);
	not 	XG3672 	(WX6782,WX7468);
	not 	XG3673 	(WX6768,WX7468);
	not 	XG3674 	(WX6754,WX7468);
	not 	XG3675 	(WX6740,WX7468);
	not 	XG3676 	(WX6726,WX7468);
	not 	XG3677 	(WX6712,WX7468);
	not 	XG3678 	(WX6698,WX7468);
	not 	XG3679 	(WX6684,WX7468);
	not 	XG3680 	(WX6670,WX7468);
	not 	XG3681 	(WX6656,WX7468);
	not 	XG3682 	(WX6642,WX7468);
	not 	XG3683 	(WX6628,WX7468);
	not 	XG3684 	(WX6614,WX7468);
	not 	XG3685 	(WX6600,WX7468);
	not 	XG3686 	(WX6586,WX7468);
	not 	XG3687 	(WX6572,WX7468);
	not 	XG3688 	(WX6558,WX7468);
	not 	XG3689 	(WX6544,WX7468);
	not 	XG3690 	(WX6530,WX7468);
	not 	XG3691 	(WX6516,WX7468);
	not 	XG3692 	(WX6502,WX7468);
	not 	XG3693 	(WX5643,WX6175);
	not 	XG3694 	(WX5629,WX6175);
	not 	XG3695 	(WX5615,WX6175);
	not 	XG3696 	(WX5601,WX6175);
	not 	XG3697 	(WX5587,WX6175);
	not 	XG3698 	(WX5573,WX6175);
	not 	XG3699 	(WX5559,WX6175);
	not 	XG3700 	(WX5545,WX6175);
	not 	XG3701 	(WX5531,WX6175);
	not 	XG3702 	(WX5517,WX6175);
	not 	XG3703 	(WX5503,WX6175);
	not 	XG3704 	(WX5489,WX6175);
	not 	XG3705 	(WX5475,WX6175);
	not 	XG3706 	(WX5461,WX6175);
	not 	XG3707 	(WX5447,WX6175);
	not 	XG3708 	(WX5433,WX6175);
	not 	XG3709 	(WX5419,WX6175);
	not 	XG3710 	(WX5405,WX6175);
	not 	XG3711 	(WX5391,WX6175);
	not 	XG3712 	(WX5377,WX6175);
	not 	XG3713 	(WX5363,WX6175);
	not 	XG3714 	(WX5349,WX6175);
	not 	XG3715 	(WX5335,WX6175);
	not 	XG3716 	(WX5321,WX6175);
	not 	XG3717 	(WX5307,WX6175);
	not 	XG3718 	(WX5293,WX6175);
	not 	XG3719 	(WX5279,WX6175);
	not 	XG3720 	(WX5265,WX6175);
	not 	XG3721 	(WX5251,WX6175);
	not 	XG3722 	(WX5237,WX6175);
	not 	XG3723 	(WX5223,WX6175);
	not 	XG3724 	(WX5209,WX6175);
	not 	XG3725 	(WX4350,WX4882);
	not 	XG3726 	(WX4336,WX4882);
	not 	XG3727 	(WX4322,WX4882);
	not 	XG3728 	(WX4308,WX4882);
	not 	XG3729 	(WX4294,WX4882);
	not 	XG3730 	(WX4280,WX4882);
	not 	XG3731 	(WX4266,WX4882);
	not 	XG3732 	(WX4252,WX4882);
	not 	XG3733 	(WX4238,WX4882);
	not 	XG3734 	(WX4224,WX4882);
	not 	XG3735 	(WX4210,WX4882);
	not 	XG3736 	(WX4196,WX4882);
	not 	XG3737 	(WX4182,WX4882);
	not 	XG3738 	(WX4168,WX4882);
	not 	XG3739 	(WX4154,WX4882);
	not 	XG3740 	(WX4140,WX4882);
	not 	XG3741 	(WX4126,WX4882);
	not 	XG3742 	(WX4112,WX4882);
	not 	XG3743 	(WX4098,WX4882);
	not 	XG3744 	(WX4084,WX4882);
	not 	XG3745 	(WX4070,WX4882);
	not 	XG3746 	(WX4056,WX4882);
	not 	XG3747 	(WX4042,WX4882);
	not 	XG3748 	(WX4028,WX4882);
	not 	XG3749 	(WX4014,WX4882);
	not 	XG3750 	(WX4000,WX4882);
	not 	XG3751 	(WX3986,WX4882);
	not 	XG3752 	(WX3972,WX4882);
	not 	XG3753 	(WX3958,WX4882);
	not 	XG3754 	(WX3944,WX4882);
	not 	XG3755 	(WX3930,WX4882);
	not 	XG3756 	(WX3916,WX4882);
	not 	XG3757 	(WX3057,WX3589);
	not 	XG3758 	(WX3043,WX3589);
	not 	XG3759 	(WX3029,WX3589);
	not 	XG3760 	(WX3015,WX3589);
	not 	XG3761 	(WX3001,WX3589);
	not 	XG3762 	(WX2987,WX3589);
	not 	XG3763 	(WX2973,WX3589);
	not 	XG3764 	(WX2959,WX3589);
	not 	XG3765 	(WX2945,WX3589);
	not 	XG3766 	(WX2931,WX3589);
	not 	XG3767 	(WX2917,WX3589);
	not 	XG3768 	(WX2903,WX3589);
	not 	XG3769 	(WX2889,WX3589);
	not 	XG3770 	(WX2875,WX3589);
	not 	XG3771 	(WX2861,WX3589);
	not 	XG3772 	(WX2847,WX3589);
	not 	XG3773 	(WX2833,WX3589);
	not 	XG3774 	(WX2819,WX3589);
	not 	XG3775 	(WX2805,WX3589);
	not 	XG3776 	(WX2791,WX3589);
	not 	XG3777 	(WX2777,WX3589);
	not 	XG3778 	(WX2763,WX3589);
	not 	XG3779 	(WX2749,WX3589);
	not 	XG3780 	(WX2735,WX3589);
	not 	XG3781 	(WX2721,WX3589);
	not 	XG3782 	(WX2707,WX3589);
	not 	XG3783 	(WX2693,WX3589);
	not 	XG3784 	(WX2679,WX3589);
	not 	XG3785 	(WX2665,WX3589);
	not 	XG3786 	(WX2651,WX3589);
	not 	XG3787 	(WX2637,WX3589);
	not 	XG3788 	(WX2623,WX3589);
	not 	XG3789 	(WX1764,WX2296);
	not 	XG3790 	(WX1750,WX2296);
	not 	XG3791 	(WX1736,WX2296);
	not 	XG3792 	(WX1722,WX2296);
	not 	XG3793 	(WX1708,WX2296);
	not 	XG3794 	(WX1694,WX2296);
	not 	XG3795 	(WX1680,WX2296);
	not 	XG3796 	(WX1666,WX2296);
	not 	XG3797 	(WX1652,WX2296);
	not 	XG3798 	(WX1638,WX2296);
	not 	XG3799 	(WX1624,WX2296);
	not 	XG3800 	(WX1610,WX2296);
	not 	XG3801 	(WX1596,WX2296);
	not 	XG3802 	(WX1582,WX2296);
	not 	XG3803 	(WX1568,WX2296);
	not 	XG3804 	(WX1554,WX2296);
	not 	XG3805 	(WX1540,WX2296);
	not 	XG3806 	(WX1526,WX2296);
	not 	XG3807 	(WX1512,WX2296);
	not 	XG3808 	(WX1498,WX2296);
	not 	XG3809 	(WX1484,WX2296);
	not 	XG3810 	(WX1470,WX2296);
	not 	XG3811 	(WX1456,WX2296);
	not 	XG3812 	(WX1442,WX2296);
	not 	XG3813 	(WX1428,WX2296);
	not 	XG3814 	(WX1414,WX2296);
	not 	XG3815 	(WX1400,WX2296);
	not 	XG3816 	(WX1386,WX2296);
	not 	XG3817 	(WX1372,WX2296);
	not 	XG3818 	(WX1358,WX2296);
	not 	XG3819 	(WX1344,WX2296);
	not 	XG3820 	(WX1330,WX2296);
	not 	XG3821 	(WX471,WX1003);
	not 	XG3822 	(WX457,WX1003);
	not 	XG3823 	(WX443,WX1003);
	not 	XG3824 	(WX429,WX1003);
	not 	XG3825 	(WX415,WX1003);
	not 	XG3826 	(WX401,WX1003);
	not 	XG3827 	(WX387,WX1003);
	not 	XG3828 	(WX373,WX1003);
	not 	XG3829 	(WX359,WX1003);
	not 	XG3830 	(WX345,WX1003);
	not 	XG3831 	(WX331,WX1003);
	not 	XG3832 	(WX317,WX1003);
	not 	XG3833 	(WX303,WX1003);
	not 	XG3834 	(WX289,WX1003);
	not 	XG3835 	(WX275,WX1003);
	not 	XG3836 	(WX261,WX1003);
	not 	XG3837 	(WX247,WX1003);
	not 	XG3838 	(WX233,WX1003);
	not 	XG3839 	(WX219,WX1003);
	not 	XG3840 	(WX205,WX1003);
	not 	XG3841 	(WX191,WX1003);
	not 	XG3842 	(WX177,WX1003);
	not 	XG3843 	(WX163,WX1003);
	not 	XG3844 	(WX149,WX1003);
	not 	XG3845 	(WX135,WX1003);
	not 	XG3846 	(WX121,WX1003);
	not 	XG3847 	(WX107,WX1003);
	not 	XG3848 	(WX93,WX1003);
	not 	XG3849 	(WX79,WX1003);
	not 	XG3850 	(WX65,WX1003);
	not 	XG3851 	(WX51,WX1003);
	not 	XG3852 	(WX37,WX1003);
	not 	XG3853 	(WX10823,WX11348);
	not 	XG3854 	(WX10819,WX11348);
	not 	XG3855 	(WX10809,WX11348);
	not 	XG3856 	(WX10805,WX11348);
	not 	XG3857 	(WX10795,WX11348);
	not 	XG3858 	(WX10791,WX11348);
	not 	XG3859 	(WX10781,WX11348);
	not 	XG3860 	(WX10777,WX11348);
	not 	XG3861 	(WX10767,WX11348);
	not 	XG3862 	(WX10763,WX11348);
	not 	XG3863 	(WX10753,WX11348);
	not 	XG3864 	(WX10749,WX11348);
	not 	XG3865 	(WX10739,WX11348);
	not 	XG3866 	(WX10735,WX11348);
	not 	XG3867 	(WX10725,WX11348);
	not 	XG3868 	(WX10721,WX11348);
	not 	XG3869 	(WX10711,WX11348);
	not 	XG3870 	(WX10707,WX11348);
	not 	XG3871 	(WX10697,WX11348);
	not 	XG3872 	(WX10693,WX11348);
	not 	XG3873 	(WX10683,WX11348);
	not 	XG3874 	(WX10679,WX11348);
	not 	XG3875 	(WX10669,WX11348);
	not 	XG3876 	(WX10665,WX11348);
	not 	XG3877 	(WX10655,WX11348);
	not 	XG3878 	(WX10651,WX11348);
	not 	XG3879 	(WX10641,WX11348);
	not 	XG3880 	(WX10637,WX11348);
	not 	XG3881 	(WX10627,WX11348);
	not 	XG3882 	(WX10623,WX11348);
	not 	XG3883 	(WX10613,WX11348);
	not 	XG3884 	(WX10609,WX11348);
	not 	XG3885 	(WX10599,WX11348);
	not 	XG3886 	(WX10595,WX11348);
	not 	XG3887 	(WX10585,WX11348);
	not 	XG3888 	(WX10581,WX11348);
	not 	XG3889 	(WX10571,WX11348);
	not 	XG3890 	(WX10567,WX11348);
	not 	XG3891 	(WX10557,WX11348);
	not 	XG3892 	(WX10553,WX11348);
	not 	XG3893 	(WX10543,WX11348);
	not 	XG3894 	(WX10539,WX11348);
	not 	XG3895 	(WX10529,WX11348);
	not 	XG3896 	(WX10525,WX11348);
	not 	XG3897 	(WX10515,WX11348);
	not 	XG3898 	(WX10511,WX11348);
	not 	XG3899 	(WX10501,WX11348);
	not 	XG3900 	(WX10497,WX11348);
	not 	XG3901 	(WX10487,WX11348);
	not 	XG3902 	(WX10483,WX11348);
	not 	XG3903 	(WX10473,WX11348);
	not 	XG3904 	(WX10469,WX11348);
	not 	XG3905 	(WX10459,WX11348);
	not 	XG3906 	(WX10455,WX11348);
	not 	XG3907 	(WX10445,WX11348);
	not 	XG3908 	(WX10441,WX11348);
	not 	XG3909 	(WX10431,WX11348);
	not 	XG3910 	(WX10427,WX11348);
	not 	XG3911 	(WX10417,WX11348);
	not 	XG3912 	(WX10413,WX11348);
	not 	XG3913 	(WX10403,WX11348);
	not 	XG3914 	(WX10399,WX11348);
	not 	XG3915 	(WX10389,WX11348);
	not 	XG3916 	(WX10385,WX11348);
	not 	XG3917 	(WX11570,WX11349);
	not 	XG3918 	(WX11563,WX11349);
	not 	XG3919 	(WX11556,WX11349);
	not 	XG3920 	(WX11549,WX11349);
	not 	XG3921 	(WX11542,WX11349);
	not 	XG3922 	(WX11535,WX11349);
	not 	XG3923 	(WX11528,WX11349);
	not 	XG3924 	(WX11521,WX11349);
	not 	XG3925 	(WX11514,WX11349);
	not 	XG3926 	(WX11507,WX11349);
	not 	XG3927 	(WX11500,WX11349);
	not 	XG3928 	(WX11493,WX11349);
	not 	XG3929 	(WX11486,WX11349);
	not 	XG3930 	(WX11479,WX11349);
	not 	XG3931 	(WX11472,WX11349);
	not 	XG3932 	(WX11465,WX11349);
	not 	XG3933 	(WX11458,WX11349);
	not 	XG3934 	(WX11451,WX11349);
	not 	XG3935 	(WX11444,WX11349);
	not 	XG3936 	(WX11437,WX11349);
	not 	XG3937 	(WX11430,WX11349);
	not 	XG3938 	(WX11423,WX11349);
	not 	XG3939 	(WX11416,WX11349);
	not 	XG3940 	(WX11409,WX11349);
	not 	XG3941 	(WX11402,WX11349);
	not 	XG3942 	(WX11395,WX11349);
	not 	XG3943 	(WX11388,WX11349);
	not 	XG3944 	(WX11381,WX11349);
	not 	XG3945 	(WX11374,WX11349);
	not 	XG3946 	(WX11367,WX11349);
	not 	XG3947 	(WX11360,WX11349);
	not 	XG3948 	(WX11353,WX11349);
	not 	XG3949 	(WX9530,WX10055);
	not 	XG3950 	(WX9526,WX10055);
	not 	XG3951 	(WX9516,WX10055);
	not 	XG3952 	(WX9512,WX10055);
	not 	XG3953 	(WX9502,WX10055);
	not 	XG3954 	(WX9498,WX10055);
	not 	XG3955 	(WX9488,WX10055);
	not 	XG3956 	(WX9484,WX10055);
	not 	XG3957 	(WX9474,WX10055);
	not 	XG3958 	(WX9470,WX10055);
	not 	XG3959 	(WX9460,WX10055);
	not 	XG3960 	(WX9456,WX10055);
	not 	XG3961 	(WX9446,WX10055);
	not 	XG3962 	(WX9442,WX10055);
	not 	XG3963 	(WX9432,WX10055);
	not 	XG3964 	(WX9428,WX10055);
	not 	XG3965 	(WX9418,WX10055);
	not 	XG3966 	(WX9414,WX10055);
	not 	XG3967 	(WX9404,WX10055);
	not 	XG3968 	(WX9400,WX10055);
	not 	XG3969 	(WX9390,WX10055);
	not 	XG3970 	(WX9386,WX10055);
	not 	XG3971 	(WX9376,WX10055);
	not 	XG3972 	(WX9372,WX10055);
	not 	XG3973 	(WX9362,WX10055);
	not 	XG3974 	(WX9358,WX10055);
	not 	XG3975 	(WX9348,WX10055);
	not 	XG3976 	(WX9344,WX10055);
	not 	XG3977 	(WX9334,WX10055);
	not 	XG3978 	(WX9330,WX10055);
	not 	XG3979 	(WX9320,WX10055);
	not 	XG3980 	(WX9316,WX10055);
	not 	XG3981 	(WX9306,WX10055);
	not 	XG3982 	(WX9302,WX10055);
	not 	XG3983 	(WX9292,WX10055);
	not 	XG3984 	(WX9288,WX10055);
	not 	XG3985 	(WX9278,WX10055);
	not 	XG3986 	(WX9274,WX10055);
	not 	XG3987 	(WX9264,WX10055);
	not 	XG3988 	(WX9260,WX10055);
	not 	XG3989 	(WX9250,WX10055);
	not 	XG3990 	(WX9246,WX10055);
	not 	XG3991 	(WX9236,WX10055);
	not 	XG3992 	(WX9232,WX10055);
	not 	XG3993 	(WX9222,WX10055);
	not 	XG3994 	(WX9218,WX10055);
	not 	XG3995 	(WX9208,WX10055);
	not 	XG3996 	(WX9204,WX10055);
	not 	XG3997 	(WX9194,WX10055);
	not 	XG3998 	(WX9190,WX10055);
	not 	XG3999 	(WX9180,WX10055);
	not 	XG4000 	(WX9176,WX10055);
	not 	XG4001 	(WX9166,WX10055);
	not 	XG4002 	(WX9162,WX10055);
	not 	XG4003 	(WX9152,WX10055);
	not 	XG4004 	(WX9148,WX10055);
	not 	XG4005 	(WX9138,WX10055);
	not 	XG4006 	(WX9134,WX10055);
	not 	XG4007 	(WX9124,WX10055);
	not 	XG4008 	(WX9120,WX10055);
	not 	XG4009 	(WX9110,WX10055);
	not 	XG4010 	(WX9106,WX10055);
	not 	XG4011 	(WX9096,WX10055);
	not 	XG4012 	(WX9092,WX10055);
	not 	XG4013 	(WX10277,WX10056);
	not 	XG4014 	(WX10270,WX10056);
	not 	XG4015 	(WX10263,WX10056);
	not 	XG4016 	(WX10256,WX10056);
	not 	XG4017 	(WX10249,WX10056);
	not 	XG4018 	(WX10242,WX10056);
	not 	XG4019 	(WX10235,WX10056);
	not 	XG4020 	(WX10228,WX10056);
	not 	XG4021 	(WX10221,WX10056);
	not 	XG4022 	(WX10214,WX10056);
	not 	XG4023 	(WX10207,WX10056);
	not 	XG4024 	(WX10200,WX10056);
	not 	XG4025 	(WX10193,WX10056);
	not 	XG4026 	(WX10186,WX10056);
	not 	XG4027 	(WX10179,WX10056);
	not 	XG4028 	(WX10172,WX10056);
	not 	XG4029 	(WX10165,WX10056);
	not 	XG4030 	(WX10158,WX10056);
	not 	XG4031 	(WX10151,WX10056);
	not 	XG4032 	(WX10144,WX10056);
	not 	XG4033 	(WX10137,WX10056);
	not 	XG4034 	(WX10130,WX10056);
	not 	XG4035 	(WX10123,WX10056);
	not 	XG4036 	(WX10116,WX10056);
	not 	XG4037 	(WX10109,WX10056);
	not 	XG4038 	(WX10102,WX10056);
	not 	XG4039 	(WX10095,WX10056);
	not 	XG4040 	(WX10088,WX10056);
	not 	XG4041 	(WX10081,WX10056);
	not 	XG4042 	(WX10074,WX10056);
	not 	XG4043 	(WX10067,WX10056);
	not 	XG4044 	(WX10060,WX10056);
	not 	XG4045 	(WX8237,WX8762);
	not 	XG4046 	(WX8233,WX8762);
	not 	XG4047 	(WX8223,WX8762);
	not 	XG4048 	(WX8219,WX8762);
	not 	XG4049 	(WX8209,WX8762);
	not 	XG4050 	(WX8205,WX8762);
	not 	XG4051 	(WX8195,WX8762);
	not 	XG4052 	(WX8191,WX8762);
	not 	XG4053 	(WX8181,WX8762);
	not 	XG4054 	(WX8177,WX8762);
	not 	XG4055 	(WX8167,WX8762);
	not 	XG4056 	(WX8163,WX8762);
	not 	XG4057 	(WX8153,WX8762);
	not 	XG4058 	(WX8149,WX8762);
	not 	XG4059 	(WX8139,WX8762);
	not 	XG4060 	(WX8135,WX8762);
	not 	XG4061 	(WX8125,WX8762);
	not 	XG4062 	(WX8121,WX8762);
	not 	XG4063 	(WX8111,WX8762);
	not 	XG4064 	(WX8107,WX8762);
	not 	XG4065 	(WX8097,WX8762);
	not 	XG4066 	(WX8093,WX8762);
	not 	XG4067 	(WX8083,WX8762);
	not 	XG4068 	(WX8079,WX8762);
	not 	XG4069 	(WX8069,WX8762);
	not 	XG4070 	(WX8065,WX8762);
	not 	XG4071 	(WX8055,WX8762);
	not 	XG4072 	(WX8051,WX8762);
	not 	XG4073 	(WX8041,WX8762);
	not 	XG4074 	(WX8037,WX8762);
	not 	XG4075 	(WX8027,WX8762);
	not 	XG4076 	(WX8023,WX8762);
	not 	XG4077 	(WX8013,WX8762);
	not 	XG4078 	(WX8009,WX8762);
	not 	XG4079 	(WX7999,WX8762);
	not 	XG4080 	(WX7995,WX8762);
	not 	XG4081 	(WX7985,WX8762);
	not 	XG4082 	(WX7981,WX8762);
	not 	XG4083 	(WX7971,WX8762);
	not 	XG4084 	(WX7967,WX8762);
	not 	XG4085 	(WX7957,WX8762);
	not 	XG4086 	(WX7953,WX8762);
	not 	XG4087 	(WX7943,WX8762);
	not 	XG4088 	(WX7939,WX8762);
	not 	XG4089 	(WX7929,WX8762);
	not 	XG4090 	(WX7925,WX8762);
	not 	XG4091 	(WX7915,WX8762);
	not 	XG4092 	(WX7911,WX8762);
	not 	XG4093 	(WX7901,WX8762);
	not 	XG4094 	(WX7897,WX8762);
	not 	XG4095 	(WX7887,WX8762);
	not 	XG4096 	(WX7883,WX8762);
	not 	XG4097 	(WX7873,WX8762);
	not 	XG4098 	(WX7869,WX8762);
	not 	XG4099 	(WX7859,WX8762);
	not 	XG4100 	(WX7855,WX8762);
	not 	XG4101 	(WX7845,WX8762);
	not 	XG4102 	(WX7841,WX8762);
	not 	XG4103 	(WX7831,WX8762);
	not 	XG4104 	(WX7827,WX8762);
	not 	XG4105 	(WX7817,WX8762);
	not 	XG4106 	(WX7813,WX8762);
	not 	XG4107 	(WX7803,WX8762);
	not 	XG4108 	(WX7799,WX8762);
	not 	XG4109 	(WX8984,WX8763);
	not 	XG4110 	(WX8977,WX8763);
	not 	XG4111 	(WX8970,WX8763);
	not 	XG4112 	(WX8963,WX8763);
	not 	XG4113 	(WX8956,WX8763);
	not 	XG4114 	(WX8949,WX8763);
	not 	XG4115 	(WX8942,WX8763);
	not 	XG4116 	(WX8935,WX8763);
	not 	XG4117 	(WX8928,WX8763);
	not 	XG4118 	(WX8921,WX8763);
	not 	XG4119 	(WX8914,WX8763);
	not 	XG4120 	(WX8907,WX8763);
	not 	XG4121 	(WX8900,WX8763);
	not 	XG4122 	(WX8893,WX8763);
	not 	XG4123 	(WX8886,WX8763);
	not 	XG4124 	(WX8879,WX8763);
	not 	XG4125 	(WX8872,WX8763);
	not 	XG4126 	(WX8865,WX8763);
	not 	XG4127 	(WX8858,WX8763);
	not 	XG4128 	(WX8851,WX8763);
	not 	XG4129 	(WX8844,WX8763);
	not 	XG4130 	(WX8837,WX8763);
	not 	XG4131 	(WX8830,WX8763);
	not 	XG4132 	(WX8823,WX8763);
	not 	XG4133 	(WX8816,WX8763);
	not 	XG4134 	(WX8809,WX8763);
	not 	XG4135 	(WX8802,WX8763);
	not 	XG4136 	(WX8795,WX8763);
	not 	XG4137 	(WX8788,WX8763);
	not 	XG4138 	(WX8781,WX8763);
	not 	XG4139 	(WX8774,WX8763);
	not 	XG4140 	(WX8767,WX8763);
	not 	XG4141 	(WX6944,WX7469);
	not 	XG4142 	(WX6940,WX7469);
	not 	XG4143 	(WX6930,WX7469);
	not 	XG4144 	(WX6926,WX7469);
	not 	XG4145 	(WX6916,WX7469);
	not 	XG4146 	(WX6912,WX7469);
	not 	XG4147 	(WX6902,WX7469);
	not 	XG4148 	(WX6898,WX7469);
	not 	XG4149 	(WX6888,WX7469);
	not 	XG4150 	(WX6884,WX7469);
	not 	XG4151 	(WX6874,WX7469);
	not 	XG4152 	(WX6870,WX7469);
	not 	XG4153 	(WX6860,WX7469);
	not 	XG4154 	(WX6856,WX7469);
	not 	XG4155 	(WX6846,WX7469);
	not 	XG4156 	(WX6842,WX7469);
	not 	XG4157 	(WX6832,WX7469);
	not 	XG4158 	(WX6828,WX7469);
	not 	XG4159 	(WX6818,WX7469);
	not 	XG4160 	(WX6814,WX7469);
	not 	XG4161 	(WX6804,WX7469);
	not 	XG4162 	(WX6800,WX7469);
	not 	XG4163 	(WX6790,WX7469);
	not 	XG4164 	(WX6786,WX7469);
	not 	XG4165 	(WX6776,WX7469);
	not 	XG4166 	(WX6772,WX7469);
	not 	XG4167 	(WX6762,WX7469);
	not 	XG4168 	(WX6758,WX7469);
	not 	XG4169 	(WX6748,WX7469);
	not 	XG4170 	(WX6744,WX7469);
	not 	XG4171 	(WX6734,WX7469);
	not 	XG4172 	(WX6730,WX7469);
	not 	XG4173 	(WX6720,WX7469);
	not 	XG4174 	(WX6716,WX7469);
	not 	XG4175 	(WX6706,WX7469);
	not 	XG4176 	(WX6702,WX7469);
	not 	XG4177 	(WX6692,WX7469);
	not 	XG4178 	(WX6688,WX7469);
	not 	XG4179 	(WX6678,WX7469);
	not 	XG4180 	(WX6674,WX7469);
	not 	XG4181 	(WX6664,WX7469);
	not 	XG4182 	(WX6660,WX7469);
	not 	XG4183 	(WX6650,WX7469);
	not 	XG4184 	(WX6646,WX7469);
	not 	XG4185 	(WX6636,WX7469);
	not 	XG4186 	(WX6632,WX7469);
	not 	XG4187 	(WX6622,WX7469);
	not 	XG4188 	(WX6618,WX7469);
	not 	XG4189 	(WX6608,WX7469);
	not 	XG4190 	(WX6604,WX7469);
	not 	XG4191 	(WX6594,WX7469);
	not 	XG4192 	(WX6590,WX7469);
	not 	XG4193 	(WX6580,WX7469);
	not 	XG4194 	(WX6576,WX7469);
	not 	XG4195 	(WX6566,WX7469);
	not 	XG4196 	(WX6562,WX7469);
	not 	XG4197 	(WX6552,WX7469);
	not 	XG4198 	(WX6548,WX7469);
	not 	XG4199 	(WX6538,WX7469);
	not 	XG4200 	(WX6534,WX7469);
	not 	XG4201 	(WX6524,WX7469);
	not 	XG4202 	(WX6520,WX7469);
	not 	XG4203 	(WX6510,WX7469);
	not 	XG4204 	(WX6506,WX7469);
	not 	XG4205 	(WX7691,WX7470);
	not 	XG4206 	(WX7684,WX7470);
	not 	XG4207 	(WX7677,WX7470);
	not 	XG4208 	(WX7670,WX7470);
	not 	XG4209 	(WX7663,WX7470);
	not 	XG4210 	(WX7656,WX7470);
	not 	XG4211 	(WX7649,WX7470);
	not 	XG4212 	(WX7642,WX7470);
	not 	XG4213 	(WX7635,WX7470);
	not 	XG4214 	(WX7628,WX7470);
	not 	XG4215 	(WX7621,WX7470);
	not 	XG4216 	(WX7614,WX7470);
	not 	XG4217 	(WX7607,WX7470);
	not 	XG4218 	(WX7600,WX7470);
	not 	XG4219 	(WX7593,WX7470);
	not 	XG4220 	(WX7586,WX7470);
	not 	XG4221 	(WX7579,WX7470);
	not 	XG4222 	(WX7572,WX7470);
	not 	XG4223 	(WX7565,WX7470);
	not 	XG4224 	(WX7558,WX7470);
	not 	XG4225 	(WX7551,WX7470);
	not 	XG4226 	(WX7544,WX7470);
	not 	XG4227 	(WX7537,WX7470);
	not 	XG4228 	(WX7530,WX7470);
	not 	XG4229 	(WX7523,WX7470);
	not 	XG4230 	(WX7516,WX7470);
	not 	XG4231 	(WX7509,WX7470);
	not 	XG4232 	(WX7502,WX7470);
	not 	XG4233 	(WX7495,WX7470);
	not 	XG4234 	(WX7488,WX7470);
	not 	XG4235 	(WX7481,WX7470);
	not 	XG4236 	(WX7474,WX7470);
	not 	XG4237 	(WX5651,WX6176);
	not 	XG4238 	(WX5647,WX6176);
	not 	XG4239 	(WX5637,WX6176);
	not 	XG4240 	(WX5633,WX6176);
	not 	XG4241 	(WX5623,WX6176);
	not 	XG4242 	(WX5619,WX6176);
	not 	XG4243 	(WX5609,WX6176);
	not 	XG4244 	(WX5605,WX6176);
	not 	XG4245 	(WX5595,WX6176);
	not 	XG4246 	(WX5591,WX6176);
	not 	XG4247 	(WX5581,WX6176);
	not 	XG4248 	(WX5577,WX6176);
	not 	XG4249 	(WX5567,WX6176);
	not 	XG4250 	(WX5563,WX6176);
	not 	XG4251 	(WX5553,WX6176);
	not 	XG4252 	(WX5549,WX6176);
	not 	XG4253 	(WX5539,WX6176);
	not 	XG4254 	(WX5535,WX6176);
	not 	XG4255 	(WX5525,WX6176);
	not 	XG4256 	(WX5521,WX6176);
	not 	XG4257 	(WX5511,WX6176);
	not 	XG4258 	(WX5507,WX6176);
	not 	XG4259 	(WX5497,WX6176);
	not 	XG4260 	(WX5493,WX6176);
	not 	XG4261 	(WX5483,WX6176);
	not 	XG4262 	(WX5479,WX6176);
	not 	XG4263 	(WX5469,WX6176);
	not 	XG4264 	(WX5465,WX6176);
	not 	XG4265 	(WX5455,WX6176);
	not 	XG4266 	(WX5451,WX6176);
	not 	XG4267 	(WX5441,WX6176);
	not 	XG4268 	(WX5437,WX6176);
	not 	XG4269 	(WX5427,WX6176);
	not 	XG4270 	(WX5423,WX6176);
	not 	XG4271 	(WX5413,WX6176);
	not 	XG4272 	(WX5409,WX6176);
	not 	XG4273 	(WX5399,WX6176);
	not 	XG4274 	(WX5395,WX6176);
	not 	XG4275 	(WX5385,WX6176);
	not 	XG4276 	(WX5381,WX6176);
	not 	XG4277 	(WX5371,WX6176);
	not 	XG4278 	(WX5367,WX6176);
	not 	XG4279 	(WX5357,WX6176);
	not 	XG4280 	(WX5353,WX6176);
	not 	XG4281 	(WX5343,WX6176);
	not 	XG4282 	(WX5339,WX6176);
	not 	XG4283 	(WX5329,WX6176);
	not 	XG4284 	(WX5325,WX6176);
	not 	XG4285 	(WX5315,WX6176);
	not 	XG4286 	(WX5311,WX6176);
	not 	XG4287 	(WX5301,WX6176);
	not 	XG4288 	(WX5297,WX6176);
	not 	XG4289 	(WX5287,WX6176);
	not 	XG4290 	(WX5283,WX6176);
	not 	XG4291 	(WX5273,WX6176);
	not 	XG4292 	(WX5269,WX6176);
	not 	XG4293 	(WX5259,WX6176);
	not 	XG4294 	(WX5255,WX6176);
	not 	XG4295 	(WX5245,WX6176);
	not 	XG4296 	(WX5241,WX6176);
	not 	XG4297 	(WX5231,WX6176);
	not 	XG4298 	(WX5227,WX6176);
	not 	XG4299 	(WX5217,WX6176);
	not 	XG4300 	(WX5213,WX6176);
	not 	XG4301 	(WX6398,WX6177);
	not 	XG4302 	(WX6391,WX6177);
	not 	XG4303 	(WX6384,WX6177);
	not 	XG4304 	(WX6377,WX6177);
	not 	XG4305 	(WX6370,WX6177);
	not 	XG4306 	(WX6363,WX6177);
	not 	XG4307 	(WX6356,WX6177);
	not 	XG4308 	(WX6349,WX6177);
	not 	XG4309 	(WX6342,WX6177);
	not 	XG4310 	(WX6335,WX6177);
	not 	XG4311 	(WX6328,WX6177);
	not 	XG4312 	(WX6321,WX6177);
	not 	XG4313 	(WX6314,WX6177);
	not 	XG4314 	(WX6307,WX6177);
	not 	XG4315 	(WX6300,WX6177);
	not 	XG4316 	(WX6293,WX6177);
	not 	XG4317 	(WX6286,WX6177);
	not 	XG4318 	(WX6279,WX6177);
	not 	XG4319 	(WX6272,WX6177);
	not 	XG4320 	(WX6265,WX6177);
	not 	XG4321 	(WX6258,WX6177);
	not 	XG4322 	(WX6251,WX6177);
	not 	XG4323 	(WX6244,WX6177);
	not 	XG4324 	(WX6237,WX6177);
	not 	XG4325 	(WX6230,WX6177);
	not 	XG4326 	(WX6223,WX6177);
	not 	XG4327 	(WX6216,WX6177);
	not 	XG4328 	(WX6209,WX6177);
	not 	XG4329 	(WX6202,WX6177);
	not 	XG4330 	(WX6195,WX6177);
	not 	XG4331 	(WX6188,WX6177);
	not 	XG4332 	(WX6181,WX6177);
	not 	XG4333 	(WX4358,WX4883);
	not 	XG4334 	(WX4354,WX4883);
	not 	XG4335 	(WX4344,WX4883);
	not 	XG4336 	(WX4340,WX4883);
	not 	XG4337 	(WX4330,WX4883);
	not 	XG4338 	(WX4326,WX4883);
	not 	XG4339 	(WX4316,WX4883);
	not 	XG4340 	(WX4312,WX4883);
	not 	XG4341 	(WX4302,WX4883);
	not 	XG4342 	(WX4298,WX4883);
	not 	XG4343 	(WX4288,WX4883);
	not 	XG4344 	(WX4284,WX4883);
	not 	XG4345 	(WX4274,WX4883);
	not 	XG4346 	(WX4270,WX4883);
	not 	XG4347 	(WX4260,WX4883);
	not 	XG4348 	(WX4256,WX4883);
	not 	XG4349 	(WX4246,WX4883);
	not 	XG4350 	(WX4242,WX4883);
	not 	XG4351 	(WX4232,WX4883);
	not 	XG4352 	(WX4228,WX4883);
	not 	XG4353 	(WX4218,WX4883);
	not 	XG4354 	(WX4214,WX4883);
	not 	XG4355 	(WX4204,WX4883);
	not 	XG4356 	(WX4200,WX4883);
	not 	XG4357 	(WX4190,WX4883);
	not 	XG4358 	(WX4186,WX4883);
	not 	XG4359 	(WX4176,WX4883);
	not 	XG4360 	(WX4172,WX4883);
	not 	XG4361 	(WX4162,WX4883);
	not 	XG4362 	(WX4158,WX4883);
	not 	XG4363 	(WX4148,WX4883);
	not 	XG4364 	(WX4144,WX4883);
	not 	XG4365 	(WX4134,WX4883);
	not 	XG4366 	(WX4130,WX4883);
	not 	XG4367 	(WX4120,WX4883);
	not 	XG4368 	(WX4116,WX4883);
	not 	XG4369 	(WX4106,WX4883);
	not 	XG4370 	(WX4102,WX4883);
	not 	XG4371 	(WX4092,WX4883);
	not 	XG4372 	(WX4088,WX4883);
	not 	XG4373 	(WX4078,WX4883);
	not 	XG4374 	(WX4074,WX4883);
	not 	XG4375 	(WX4064,WX4883);
	not 	XG4376 	(WX4060,WX4883);
	not 	XG4377 	(WX4050,WX4883);
	not 	XG4378 	(WX4046,WX4883);
	not 	XG4379 	(WX4036,WX4883);
	not 	XG4380 	(WX4032,WX4883);
	not 	XG4381 	(WX4022,WX4883);
	not 	XG4382 	(WX4018,WX4883);
	not 	XG4383 	(WX4008,WX4883);
	not 	XG4384 	(WX4004,WX4883);
	not 	XG4385 	(WX3994,WX4883);
	not 	XG4386 	(WX3990,WX4883);
	not 	XG4387 	(WX3980,WX4883);
	not 	XG4388 	(WX3976,WX4883);
	not 	XG4389 	(WX3966,WX4883);
	not 	XG4390 	(WX3962,WX4883);
	not 	XG4391 	(WX3952,WX4883);
	not 	XG4392 	(WX3948,WX4883);
	not 	XG4393 	(WX3938,WX4883);
	not 	XG4394 	(WX3934,WX4883);
	not 	XG4395 	(WX3924,WX4883);
	not 	XG4396 	(WX3920,WX4883);
	not 	XG4397 	(WX5105,WX4884);
	not 	XG4398 	(WX5098,WX4884);
	not 	XG4399 	(WX5091,WX4884);
	not 	XG4400 	(WX5084,WX4884);
	not 	XG4401 	(WX5077,WX4884);
	not 	XG4402 	(WX5070,WX4884);
	not 	XG4403 	(WX5063,WX4884);
	not 	XG4404 	(WX5056,WX4884);
	not 	XG4405 	(WX5049,WX4884);
	not 	XG4406 	(WX5042,WX4884);
	not 	XG4407 	(WX5035,WX4884);
	not 	XG4408 	(WX5028,WX4884);
	not 	XG4409 	(WX5021,WX4884);
	not 	XG4410 	(WX5014,WX4884);
	not 	XG4411 	(WX5007,WX4884);
	not 	XG4412 	(WX5000,WX4884);
	not 	XG4413 	(WX4993,WX4884);
	not 	XG4414 	(WX4986,WX4884);
	not 	XG4415 	(WX4979,WX4884);
	not 	XG4416 	(WX4972,WX4884);
	not 	XG4417 	(WX4965,WX4884);
	not 	XG4418 	(WX4958,WX4884);
	not 	XG4419 	(WX4951,WX4884);
	not 	XG4420 	(WX4944,WX4884);
	not 	XG4421 	(WX4937,WX4884);
	not 	XG4422 	(WX4930,WX4884);
	not 	XG4423 	(WX4923,WX4884);
	not 	XG4424 	(WX4916,WX4884);
	not 	XG4425 	(WX4909,WX4884);
	not 	XG4426 	(WX4902,WX4884);
	not 	XG4427 	(WX4895,WX4884);
	not 	XG4428 	(WX4888,WX4884);
	not 	XG4429 	(WX3065,WX3590);
	not 	XG4430 	(WX3061,WX3590);
	not 	XG4431 	(WX3051,WX3590);
	not 	XG4432 	(WX3047,WX3590);
	not 	XG4433 	(WX3037,WX3590);
	not 	XG4434 	(WX3033,WX3590);
	not 	XG4435 	(WX3023,WX3590);
	not 	XG4436 	(WX3019,WX3590);
	not 	XG4437 	(WX3009,WX3590);
	not 	XG4438 	(WX3005,WX3590);
	not 	XG4439 	(WX2995,WX3590);
	not 	XG4440 	(WX2991,WX3590);
	not 	XG4441 	(WX2981,WX3590);
	not 	XG4442 	(WX2977,WX3590);
	not 	XG4443 	(WX2967,WX3590);
	not 	XG4444 	(WX2963,WX3590);
	not 	XG4445 	(WX2953,WX3590);
	not 	XG4446 	(WX2949,WX3590);
	not 	XG4447 	(WX2939,WX3590);
	not 	XG4448 	(WX2935,WX3590);
	not 	XG4449 	(WX2925,WX3590);
	not 	XG4450 	(WX2921,WX3590);
	not 	XG4451 	(WX2911,WX3590);
	not 	XG4452 	(WX2907,WX3590);
	not 	XG4453 	(WX2897,WX3590);
	not 	XG4454 	(WX2893,WX3590);
	not 	XG4455 	(WX2883,WX3590);
	not 	XG4456 	(WX2879,WX3590);
	not 	XG4457 	(WX2869,WX3590);
	not 	XG4458 	(WX2865,WX3590);
	not 	XG4459 	(WX2855,WX3590);
	not 	XG4460 	(WX2851,WX3590);
	not 	XG4461 	(WX2841,WX3590);
	not 	XG4462 	(WX2837,WX3590);
	not 	XG4463 	(WX2827,WX3590);
	not 	XG4464 	(WX2823,WX3590);
	not 	XG4465 	(WX2813,WX3590);
	not 	XG4466 	(WX2809,WX3590);
	not 	XG4467 	(WX2799,WX3590);
	not 	XG4468 	(WX2795,WX3590);
	not 	XG4469 	(WX2785,WX3590);
	not 	XG4470 	(WX2781,WX3590);
	not 	XG4471 	(WX2771,WX3590);
	not 	XG4472 	(WX2767,WX3590);
	not 	XG4473 	(WX2757,WX3590);
	not 	XG4474 	(WX2753,WX3590);
	not 	XG4475 	(WX2743,WX3590);
	not 	XG4476 	(WX2739,WX3590);
	not 	XG4477 	(WX2729,WX3590);
	not 	XG4478 	(WX2725,WX3590);
	not 	XG4479 	(WX2715,WX3590);
	not 	XG4480 	(WX2711,WX3590);
	not 	XG4481 	(WX2701,WX3590);
	not 	XG4482 	(WX2697,WX3590);
	not 	XG4483 	(WX2687,WX3590);
	not 	XG4484 	(WX2683,WX3590);
	not 	XG4485 	(WX2673,WX3590);
	not 	XG4486 	(WX2669,WX3590);
	not 	XG4487 	(WX2659,WX3590);
	not 	XG4488 	(WX2655,WX3590);
	not 	XG4489 	(WX2645,WX3590);
	not 	XG4490 	(WX2641,WX3590);
	not 	XG4491 	(WX2631,WX3590);
	not 	XG4492 	(WX2627,WX3590);
	not 	XG4493 	(WX3812,WX3591);
	not 	XG4494 	(WX3805,WX3591);
	not 	XG4495 	(WX3798,WX3591);
	not 	XG4496 	(WX3791,WX3591);
	not 	XG4497 	(WX3784,WX3591);
	not 	XG4498 	(WX3777,WX3591);
	not 	XG4499 	(WX3770,WX3591);
	not 	XG4500 	(WX3763,WX3591);
	not 	XG4501 	(WX3756,WX3591);
	not 	XG4502 	(WX3749,WX3591);
	not 	XG4503 	(WX3742,WX3591);
	not 	XG4504 	(WX3735,WX3591);
	not 	XG4505 	(WX3728,WX3591);
	not 	XG4506 	(WX3721,WX3591);
	not 	XG4507 	(WX3714,WX3591);
	not 	XG4508 	(WX3707,WX3591);
	not 	XG4509 	(WX3700,WX3591);
	not 	XG4510 	(WX3693,WX3591);
	not 	XG4511 	(WX3686,WX3591);
	not 	XG4512 	(WX3679,WX3591);
	not 	XG4513 	(WX3672,WX3591);
	not 	XG4514 	(WX3665,WX3591);
	not 	XG4515 	(WX3658,WX3591);
	not 	XG4516 	(WX3651,WX3591);
	not 	XG4517 	(WX3644,WX3591);
	not 	XG4518 	(WX3637,WX3591);
	not 	XG4519 	(WX3630,WX3591);
	not 	XG4520 	(WX3623,WX3591);
	not 	XG4521 	(WX3616,WX3591);
	not 	XG4522 	(WX3609,WX3591);
	not 	XG4523 	(WX3602,WX3591);
	not 	XG4524 	(WX3595,WX3591);
	not 	XG4525 	(WX1772,WX2297);
	not 	XG4526 	(WX1768,WX2297);
	not 	XG4527 	(WX1758,WX2297);
	not 	XG4528 	(WX1754,WX2297);
	not 	XG4529 	(WX1744,WX2297);
	not 	XG4530 	(WX1740,WX2297);
	not 	XG4531 	(WX1730,WX2297);
	not 	XG4532 	(WX1726,WX2297);
	not 	XG4533 	(WX1716,WX2297);
	not 	XG4534 	(WX1712,WX2297);
	not 	XG4535 	(WX1702,WX2297);
	not 	XG4536 	(WX1698,WX2297);
	not 	XG4537 	(WX1688,WX2297);
	not 	XG4538 	(WX1684,WX2297);
	not 	XG4539 	(WX1674,WX2297);
	not 	XG4540 	(WX1670,WX2297);
	not 	XG4541 	(WX1660,WX2297);
	not 	XG4542 	(WX1656,WX2297);
	not 	XG4543 	(WX1646,WX2297);
	not 	XG4544 	(WX1642,WX2297);
	not 	XG4545 	(WX1632,WX2297);
	not 	XG4546 	(WX1628,WX2297);
	not 	XG4547 	(WX1618,WX2297);
	not 	XG4548 	(WX1614,WX2297);
	not 	XG4549 	(WX1604,WX2297);
	not 	XG4550 	(WX1600,WX2297);
	not 	XG4551 	(WX1590,WX2297);
	not 	XG4552 	(WX1586,WX2297);
	not 	XG4553 	(WX1576,WX2297);
	not 	XG4554 	(WX1572,WX2297);
	not 	XG4555 	(WX1562,WX2297);
	not 	XG4556 	(WX1558,WX2297);
	not 	XG4557 	(WX1548,WX2297);
	not 	XG4558 	(WX1544,WX2297);
	not 	XG4559 	(WX1534,WX2297);
	not 	XG4560 	(WX1530,WX2297);
	not 	XG4561 	(WX1520,WX2297);
	not 	XG4562 	(WX1516,WX2297);
	not 	XG4563 	(WX1506,WX2297);
	not 	XG4564 	(WX1502,WX2297);
	not 	XG4565 	(WX1492,WX2297);
	not 	XG4566 	(WX1488,WX2297);
	not 	XG4567 	(WX1478,WX2297);
	not 	XG4568 	(WX1474,WX2297);
	not 	XG4569 	(WX1464,WX2297);
	not 	XG4570 	(WX1460,WX2297);
	not 	XG4571 	(WX1450,WX2297);
	not 	XG4572 	(WX1446,WX2297);
	not 	XG4573 	(WX1436,WX2297);
	not 	XG4574 	(WX1432,WX2297);
	not 	XG4575 	(WX1422,WX2297);
	not 	XG4576 	(WX1418,WX2297);
	not 	XG4577 	(WX1408,WX2297);
	not 	XG4578 	(WX1404,WX2297);
	not 	XG4579 	(WX1394,WX2297);
	not 	XG4580 	(WX1390,WX2297);
	not 	XG4581 	(WX1380,WX2297);
	not 	XG4582 	(WX1376,WX2297);
	not 	XG4583 	(WX1366,WX2297);
	not 	XG4584 	(WX1362,WX2297);
	not 	XG4585 	(WX1352,WX2297);
	not 	XG4586 	(WX1348,WX2297);
	not 	XG4587 	(WX1338,WX2297);
	not 	XG4588 	(WX1334,WX2297);
	not 	XG4589 	(WX2519,WX2298);
	not 	XG4590 	(WX2512,WX2298);
	not 	XG4591 	(WX2505,WX2298);
	not 	XG4592 	(WX2498,WX2298);
	not 	XG4593 	(WX2491,WX2298);
	not 	XG4594 	(WX2484,WX2298);
	not 	XG4595 	(WX2477,WX2298);
	not 	XG4596 	(WX2470,WX2298);
	not 	XG4597 	(WX2463,WX2298);
	not 	XG4598 	(WX2456,WX2298);
	not 	XG4599 	(WX2449,WX2298);
	not 	XG4600 	(WX2442,WX2298);
	not 	XG4601 	(WX2435,WX2298);
	not 	XG4602 	(WX2428,WX2298);
	not 	XG4603 	(WX2421,WX2298);
	not 	XG4604 	(WX2414,WX2298);
	not 	XG4605 	(WX2407,WX2298);
	not 	XG4606 	(WX2400,WX2298);
	not 	XG4607 	(WX2393,WX2298);
	not 	XG4608 	(WX2386,WX2298);
	not 	XG4609 	(WX2379,WX2298);
	not 	XG4610 	(WX2372,WX2298);
	not 	XG4611 	(WX2365,WX2298);
	not 	XG4612 	(WX2358,WX2298);
	not 	XG4613 	(WX2351,WX2298);
	not 	XG4614 	(WX2344,WX2298);
	not 	XG4615 	(WX2337,WX2298);
	not 	XG4616 	(WX2330,WX2298);
	not 	XG4617 	(WX2323,WX2298);
	not 	XG4618 	(WX2316,WX2298);
	not 	XG4619 	(WX2309,WX2298);
	not 	XG4620 	(WX2302,WX2298);
	not 	XG4621 	(WX479,WX1004);
	not 	XG4622 	(WX475,WX1004);
	not 	XG4623 	(WX465,WX1004);
	not 	XG4624 	(WX461,WX1004);
	not 	XG4625 	(WX451,WX1004);
	not 	XG4626 	(WX447,WX1004);
	not 	XG4627 	(WX437,WX1004);
	not 	XG4628 	(WX433,WX1004);
	not 	XG4629 	(WX423,WX1004);
	not 	XG4630 	(WX419,WX1004);
	not 	XG4631 	(WX409,WX1004);
	not 	XG4632 	(WX405,WX1004);
	not 	XG4633 	(WX395,WX1004);
	not 	XG4634 	(WX391,WX1004);
	not 	XG4635 	(WX381,WX1004);
	not 	XG4636 	(WX377,WX1004);
	not 	XG4637 	(WX367,WX1004);
	not 	XG4638 	(WX363,WX1004);
	not 	XG4639 	(WX353,WX1004);
	not 	XG4640 	(WX349,WX1004);
	not 	XG4641 	(WX339,WX1004);
	not 	XG4642 	(WX335,WX1004);
	not 	XG4643 	(WX325,WX1004);
	not 	XG4644 	(WX321,WX1004);
	not 	XG4645 	(WX311,WX1004);
	not 	XG4646 	(WX307,WX1004);
	not 	XG4647 	(WX297,WX1004);
	not 	XG4648 	(WX293,WX1004);
	not 	XG4649 	(WX283,WX1004);
	not 	XG4650 	(WX279,WX1004);
	not 	XG4651 	(WX269,WX1004);
	not 	XG4652 	(WX265,WX1004);
	not 	XG4653 	(WX255,WX1004);
	not 	XG4654 	(WX251,WX1004);
	not 	XG4655 	(WX241,WX1004);
	not 	XG4656 	(WX237,WX1004);
	not 	XG4657 	(WX227,WX1004);
	not 	XG4658 	(WX223,WX1004);
	not 	XG4659 	(WX213,WX1004);
	not 	XG4660 	(WX209,WX1004);
	not 	XG4661 	(WX199,WX1004);
	not 	XG4662 	(WX195,WX1004);
	not 	XG4663 	(WX185,WX1004);
	not 	XG4664 	(WX181,WX1004);
	not 	XG4665 	(WX171,WX1004);
	not 	XG4666 	(WX167,WX1004);
	not 	XG4667 	(WX157,WX1004);
	not 	XG4668 	(WX153,WX1004);
	not 	XG4669 	(WX143,WX1004);
	not 	XG4670 	(WX139,WX1004);
	not 	XG4671 	(WX129,WX1004);
	not 	XG4672 	(WX125,WX1004);
	not 	XG4673 	(WX115,WX1004);
	not 	XG4674 	(WX111,WX1004);
	not 	XG4675 	(WX101,WX1004);
	not 	XG4676 	(WX97,WX1004);
	not 	XG4677 	(WX87,WX1004);
	not 	XG4678 	(WX83,WX1004);
	not 	XG4679 	(WX73,WX1004);
	not 	XG4680 	(WX69,WX1004);
	not 	XG4681 	(WX59,WX1004);
	not 	XG4682 	(WX55,WX1004);
	not 	XG4683 	(WX45,WX1004);
	not 	XG4684 	(WX41,WX1004);
	not 	XG4685 	(WX1226,WX1005);
	not 	XG4686 	(WX1219,WX1005);
	not 	XG4687 	(WX1212,WX1005);
	not 	XG4688 	(WX1205,WX1005);
	not 	XG4689 	(WX1198,WX1005);
	not 	XG4690 	(WX1191,WX1005);
	not 	XG4691 	(WX1184,WX1005);
	not 	XG4692 	(WX1177,WX1005);
	not 	XG4693 	(WX1170,WX1005);
	not 	XG4694 	(WX1163,WX1005);
	not 	XG4695 	(WX1156,WX1005);
	not 	XG4696 	(WX1149,WX1005);
	not 	XG4697 	(WX1142,WX1005);
	not 	XG4698 	(WX1135,WX1005);
	not 	XG4699 	(WX1128,WX1005);
	not 	XG4700 	(WX1121,WX1005);
	not 	XG4701 	(WX1114,WX1005);
	not 	XG4702 	(WX1107,WX1005);
	not 	XG4703 	(WX1100,WX1005);
	not 	XG4704 	(WX1093,WX1005);
	not 	XG4705 	(WX1086,WX1005);
	not 	XG4706 	(WX1079,WX1005);
	not 	XG4707 	(WX1072,WX1005);
	not 	XG4708 	(WX1065,WX1005);
	not 	XG4709 	(WX1058,WX1005);
	not 	XG4710 	(WX1051,WX1005);
	not 	XG4711 	(WX1044,WX1005);
	not 	XG4712 	(WX1037,WX1005);
	not 	XG4713 	(WX1030,WX1005);
	not 	XG4714 	(WX1023,WX1005);
	not 	XG4715 	(WX1016,WX1005);
	not 	XG4716 	(WX1009,WX1005);
	nand 	XG4717 	(II35006,II35004,WX11243);
	nand 	XG4718 	(II34975,II34973,WX11241);
	nand 	XG4719 	(II34944,II34942,WX11239);
	nand 	XG4720 	(II34913,II34911,WX11237);
	nand 	XG4721 	(II34882,II34880,WX11235);
	nand 	XG4722 	(II34851,II34849,WX11233);
	nand 	XG4723 	(II34820,II34818,WX11231);
	nand 	XG4724 	(II34789,II34787,WX11229);
	nand 	XG4725 	(II34758,II34756,WX11227);
	nand 	XG4726 	(II34727,II34725,WX11225);
	nand 	XG4727 	(II34696,II34694,WX11223);
	nand 	XG4728 	(II34665,II34663,WX11221);
	nand 	XG4729 	(II34634,II34632,WX11219);
	nand 	XG4730 	(II34603,II34601,WX11217);
	nand 	XG4731 	(II34572,II34570,WX11215);
	nand 	XG4732 	(II34541,II34539,WX11213);
	nand 	XG4733 	(II34510,II34508,WX11211);
	nand 	XG4734 	(II34479,II34477,WX11209);
	nand 	XG4735 	(II34448,II34446,WX11207);
	nand 	XG4736 	(II34417,II34415,WX11205);
	nand 	XG4737 	(II34386,II34384,WX11203);
	nand 	XG4738 	(II34355,II34353,WX11201);
	nand 	XG4739 	(II34324,II34322,WX11199);
	nand 	XG4740 	(II34293,II34291,WX11197);
	nand 	XG4741 	(II34262,II34260,WX11195);
	nand 	XG4742 	(II34231,II34229,WX11193);
	nand 	XG4743 	(II34200,II34198,WX11191);
	nand 	XG4744 	(II34169,II34167,WX11189);
	nand 	XG4745 	(II34138,II34136,WX11187);
	nand 	XG4746 	(II34107,II34105,WX11185);
	nand 	XG4747 	(II34076,II34074,WX11183);
	nand 	XG4748 	(II34045,II34043,WX11181);
	nand 	XG4749 	(II34989,WX11051,WX11346);
	nand 	XG4750 	(II34958,WX11049,WX11346);
	nand 	XG4751 	(II34927,WX11047,WX11346);
	nand 	XG4752 	(II34896,WX11045,WX11346);
	nand 	XG4753 	(II34865,WX11043,WX11346);
	nand 	XG4754 	(II34834,WX11041,WX11346);
	nand 	XG4755 	(II34803,WX11039,WX11346);
	nand 	XG4756 	(II34772,WX11037,WX11346);
	nand 	XG4757 	(II34741,WX11035,WX11346);
	nand 	XG4758 	(II34710,WX11033,WX11346);
	nand 	XG4759 	(II34679,WX11031,WX11346);
	nand 	XG4760 	(II34648,WX11029,WX11346);
	nand 	XG4761 	(II34617,WX11027,WX11346);
	nand 	XG4762 	(II34586,WX11025,WX11346);
	nand 	XG4763 	(II34555,WX11023,WX11346);
	nand 	XG4764 	(II34524,WX11021,WX11346);
	nand 	XG4765 	(II34493,WX11019,WX11345);
	nand 	XG4766 	(II34462,WX11017,WX11345);
	nand 	XG4767 	(II34431,WX11015,WX11345);
	nand 	XG4768 	(II34400,WX11013,WX11345);
	nand 	XG4769 	(II34369,WX11011,WX11345);
	nand 	XG4770 	(II34338,WX11009,WX11345);
	nand 	XG4771 	(II34307,WX11007,WX11345);
	nand 	XG4772 	(II34276,WX11005,WX11345);
	nand 	XG4773 	(II34245,WX11003,WX11345);
	nand 	XG4774 	(II34214,WX11001,WX11345);
	nand 	XG4775 	(II34183,WX10999,WX11345);
	nand 	XG4776 	(II34152,WX10997,WX11345);
	nand 	XG4777 	(II34121,WX10995,WX11345);
	nand 	XG4778 	(II34090,WX10993,WX11345);
	nand 	XG4779 	(II34059,WX10991,WX11345);
	nand 	XG4780 	(II34028,WX10989,WX11345);
	and 	XG4781 	(WX10821,WX11348,WX10891);
	and 	XG4782 	(WX10807,WX11348,WX10889);
	and 	XG4783 	(WX10793,WX11348,WX10887);
	and 	XG4784 	(WX10779,WX11348,WX10885);
	and 	XG4785 	(WX10765,WX11348,WX10883);
	and 	XG4786 	(WX10751,WX11348,WX10881);
	and 	XG4787 	(WX10737,WX11348,WX10879);
	and 	XG4788 	(WX10723,WX11348,WX10877);
	and 	XG4789 	(WX10709,WX11348,WX10875);
	and 	XG4790 	(WX10695,WX11348,WX10873);
	and 	XG4791 	(WX10681,WX11348,WX10871);
	and 	XG4792 	(WX10667,WX11348,WX10869);
	and 	XG4793 	(WX10653,WX11348,WX10867);
	and 	XG4794 	(WX10639,WX11348,WX10865);
	and 	XG4795 	(WX10625,WX11348,WX10863);
	and 	XG4796 	(WX10611,WX11348,WX10861);
	and 	XG4797 	(WX10597,WX11348,WX10859);
	and 	XG4798 	(WX10583,WX11348,WX10857);
	and 	XG4799 	(WX10569,WX11348,WX10855);
	and 	XG4800 	(WX10555,WX11348,WX10853);
	and 	XG4801 	(WX10541,WX11348,WX10851);
	and 	XG4802 	(WX10527,WX11348,WX10849);
	and 	XG4803 	(WX10513,WX11348,WX10847);
	and 	XG4804 	(WX10499,WX11348,WX10845);
	and 	XG4805 	(WX10485,WX11348,WX10843);
	and 	XG4806 	(WX10471,WX11348,WX10841);
	and 	XG4807 	(WX10457,WX11348,WX10839);
	and 	XG4808 	(WX10443,WX11348,WX10837);
	and 	XG4809 	(WX10429,WX11348,WX10835);
	and 	XG4810 	(WX10415,WX11348,WX10833);
	and 	XG4811 	(WX10401,WX11348,WX10831);
	and 	XG4812 	(WX10387,WX11348,WX10829);
	nand 	XG4813 	(II31001,II30999,WX9950);
	nand 	XG4814 	(II30970,II30968,WX9948);
	nand 	XG4815 	(II30939,II30937,WX9946);
	nand 	XG4816 	(II30908,II30906,WX9944);
	nand 	XG4817 	(II30877,II30875,WX9942);
	nand 	XG4818 	(II30846,II30844,WX9940);
	nand 	XG4819 	(II30815,II30813,WX9938);
	nand 	XG4820 	(II30784,II30782,WX9936);
	nand 	XG4821 	(II30753,II30751,WX9934);
	nand 	XG4822 	(II30722,II30720,WX9932);
	nand 	XG4823 	(II30691,II30689,WX9930);
	nand 	XG4824 	(II30660,II30658,WX9928);
	nand 	XG4825 	(II30629,II30627,WX9926);
	nand 	XG4826 	(II30598,II30596,WX9924);
	nand 	XG4827 	(II30567,II30565,WX9922);
	nand 	XG4828 	(II30536,II30534,WX9920);
	nand 	XG4829 	(II30505,II30503,WX9918);
	nand 	XG4830 	(II30474,II30472,WX9916);
	nand 	XG4831 	(II30443,II30441,WX9914);
	nand 	XG4832 	(II30412,II30410,WX9912);
	nand 	XG4833 	(II30381,II30379,WX9910);
	nand 	XG4834 	(II30350,II30348,WX9908);
	nand 	XG4835 	(II30319,II30317,WX9906);
	nand 	XG4836 	(II30288,II30286,WX9904);
	nand 	XG4837 	(II30257,II30255,WX9902);
	nand 	XG4838 	(II30226,II30224,WX9900);
	nand 	XG4839 	(II30195,II30193,WX9898);
	nand 	XG4840 	(II30164,II30162,WX9896);
	nand 	XG4841 	(II30133,II30131,WX9894);
	nand 	XG4842 	(II30102,II30100,WX9892);
	nand 	XG4843 	(II30071,II30069,WX9890);
	nand 	XG4844 	(II30040,II30038,WX9888);
	nand 	XG4845 	(II30984,WX9758,WX10053);
	nand 	XG4846 	(II30953,WX9756,WX10053);
	nand 	XG4847 	(II30922,WX9754,WX10053);
	nand 	XG4848 	(II30891,WX9752,WX10053);
	nand 	XG4849 	(II30860,WX9750,WX10053);
	nand 	XG4850 	(II30829,WX9748,WX10053);
	nand 	XG4851 	(II30798,WX9746,WX10053);
	nand 	XG4852 	(II30767,WX9744,WX10053);
	nand 	XG4853 	(II30736,WX9742,WX10053);
	nand 	XG4854 	(II30705,WX9740,WX10053);
	nand 	XG4855 	(II30674,WX9738,WX10053);
	nand 	XG4856 	(II30643,WX9736,WX10053);
	nand 	XG4857 	(II30612,WX9734,WX10053);
	nand 	XG4858 	(II30581,WX9732,WX10053);
	nand 	XG4859 	(II30550,WX9730,WX10053);
	nand 	XG4860 	(II30519,WX9728,WX10053);
	nand 	XG4861 	(II30488,WX9726,WX10052);
	nand 	XG4862 	(II30457,WX9724,WX10052);
	nand 	XG4863 	(II30426,WX9722,WX10052);
	nand 	XG4864 	(II30395,WX9720,WX10052);
	nand 	XG4865 	(II30364,WX9718,WX10052);
	nand 	XG4866 	(II30333,WX9716,WX10052);
	nand 	XG4867 	(II30302,WX9714,WX10052);
	nand 	XG4868 	(II30271,WX9712,WX10052);
	nand 	XG4869 	(II30240,WX9710,WX10052);
	nand 	XG4870 	(II30209,WX9708,WX10052);
	nand 	XG4871 	(II30178,WX9706,WX10052);
	nand 	XG4872 	(II30147,WX9704,WX10052);
	nand 	XG4873 	(II30116,WX9702,WX10052);
	nand 	XG4874 	(II30085,WX9700,WX10052);
	nand 	XG4875 	(II30054,WX9698,WX10052);
	nand 	XG4876 	(II30023,WX9696,WX10052);
	and 	XG4877 	(WX9528,WX10055,WX9598);
	and 	XG4878 	(WX9514,WX10055,WX9596);
	and 	XG4879 	(WX9500,WX10055,WX9594);
	and 	XG4880 	(WX9486,WX10055,WX9592);
	and 	XG4881 	(WX9472,WX10055,WX9590);
	and 	XG4882 	(WX9458,WX10055,WX9588);
	and 	XG4883 	(WX9444,WX10055,WX9586);
	and 	XG4884 	(WX9430,WX10055,WX9584);
	and 	XG4885 	(WX9416,WX10055,WX9582);
	and 	XG4886 	(WX9402,WX10055,WX9580);
	and 	XG4887 	(WX9388,WX10055,WX9578);
	and 	XG4888 	(WX9374,WX10055,WX9576);
	and 	XG4889 	(WX9360,WX10055,WX9574);
	and 	XG4890 	(WX9346,WX10055,WX9572);
	and 	XG4891 	(WX9332,WX10055,WX9570);
	and 	XG4892 	(WX9318,WX10055,WX9568);
	and 	XG4893 	(WX9304,WX10055,WX9566);
	and 	XG4894 	(WX9290,WX10055,WX9564);
	and 	XG4895 	(WX9276,WX10055,WX9562);
	and 	XG4896 	(WX9262,WX10055,WX9560);
	and 	XG4897 	(WX9248,WX10055,WX9558);
	and 	XG4898 	(WX9234,WX10055,WX9556);
	and 	XG4899 	(WX9220,WX10055,WX9554);
	and 	XG4900 	(WX9206,WX10055,WX9552);
	and 	XG4901 	(WX9192,WX10055,WX9550);
	and 	XG4902 	(WX9178,WX10055,WX9548);
	and 	XG4903 	(WX9164,WX10055,WX9546);
	and 	XG4904 	(WX9150,WX10055,WX9544);
	and 	XG4905 	(WX9136,WX10055,WX9542);
	and 	XG4906 	(WX9122,WX10055,WX9540);
	and 	XG4907 	(WX9108,WX10055,WX9538);
	and 	XG4908 	(WX9094,WX10055,WX9536);
	nand 	XG4909 	(II26996,II26994,WX8657);
	nand 	XG4910 	(II26965,II26963,WX8655);
	nand 	XG4911 	(II26934,II26932,WX8653);
	nand 	XG4912 	(II26903,II26901,WX8651);
	nand 	XG4913 	(II26872,II26870,WX8649);
	nand 	XG4914 	(II26841,II26839,WX8647);
	nand 	XG4915 	(II26810,II26808,WX8645);
	nand 	XG4916 	(II26779,II26777,WX8643);
	nand 	XG4917 	(II26748,II26746,WX8641);
	nand 	XG4918 	(II26717,II26715,WX8639);
	nand 	XG4919 	(II26686,II26684,WX8637);
	nand 	XG4920 	(II26655,II26653,WX8635);
	nand 	XG4921 	(II26624,II26622,WX8633);
	nand 	XG4922 	(II26593,II26591,WX8631);
	nand 	XG4923 	(II26562,II26560,WX8629);
	nand 	XG4924 	(II26531,II26529,WX8627);
	nand 	XG4925 	(II26500,II26498,WX8625);
	nand 	XG4926 	(II26469,II26467,WX8623);
	nand 	XG4927 	(II26438,II26436,WX8621);
	nand 	XG4928 	(II26407,II26405,WX8619);
	nand 	XG4929 	(II26376,II26374,WX8617);
	nand 	XG4930 	(II26345,II26343,WX8615);
	nand 	XG4931 	(II26314,II26312,WX8613);
	nand 	XG4932 	(II26283,II26281,WX8611);
	nand 	XG4933 	(II26252,II26250,WX8609);
	nand 	XG4934 	(II26221,II26219,WX8607);
	nand 	XG4935 	(II26190,II26188,WX8605);
	nand 	XG4936 	(II26159,II26157,WX8603);
	nand 	XG4937 	(II26128,II26126,WX8601);
	nand 	XG4938 	(II26097,II26095,WX8599);
	nand 	XG4939 	(II26066,II26064,WX8597);
	nand 	XG4940 	(II26035,II26033,WX8595);
	nand 	XG4941 	(II26979,WX8465,WX8760);
	nand 	XG4942 	(II26948,WX8463,WX8760);
	nand 	XG4943 	(II26917,WX8461,WX8760);
	nand 	XG4944 	(II26886,WX8459,WX8760);
	nand 	XG4945 	(II26855,WX8457,WX8760);
	nand 	XG4946 	(II26824,WX8455,WX8760);
	nand 	XG4947 	(II26793,WX8453,WX8760);
	nand 	XG4948 	(II26762,WX8451,WX8760);
	nand 	XG4949 	(II26731,WX8449,WX8760);
	nand 	XG4950 	(II26700,WX8447,WX8760);
	nand 	XG4951 	(II26669,WX8445,WX8760);
	nand 	XG4952 	(II26638,WX8443,WX8760);
	nand 	XG4953 	(II26607,WX8441,WX8760);
	nand 	XG4954 	(II26576,WX8439,WX8760);
	nand 	XG4955 	(II26545,WX8437,WX8760);
	nand 	XG4956 	(II26514,WX8435,WX8760);
	nand 	XG4957 	(II26483,WX8433,WX8759);
	nand 	XG4958 	(II26452,WX8431,WX8759);
	nand 	XG4959 	(II26421,WX8429,WX8759);
	nand 	XG4960 	(II26390,WX8427,WX8759);
	nand 	XG4961 	(II26359,WX8425,WX8759);
	nand 	XG4962 	(II26328,WX8423,WX8759);
	nand 	XG4963 	(II26297,WX8421,WX8759);
	nand 	XG4964 	(II26266,WX8419,WX8759);
	nand 	XG4965 	(II26235,WX8417,WX8759);
	nand 	XG4966 	(II26204,WX8415,WX8759);
	nand 	XG4967 	(II26173,WX8413,WX8759);
	nand 	XG4968 	(II26142,WX8411,WX8759);
	nand 	XG4969 	(II26111,WX8409,WX8759);
	nand 	XG4970 	(II26080,WX8407,WX8759);
	nand 	XG4971 	(II26049,WX8405,WX8759);
	nand 	XG4972 	(II26018,WX8403,WX8759);
	and 	XG4973 	(WX8235,WX8762,WX8305);
	and 	XG4974 	(WX8221,WX8762,WX8303);
	and 	XG4975 	(WX8207,WX8762,WX8301);
	and 	XG4976 	(WX8193,WX8762,WX8299);
	and 	XG4977 	(WX8179,WX8762,WX8297);
	and 	XG4978 	(WX8165,WX8762,WX8295);
	and 	XG4979 	(WX8151,WX8762,WX8293);
	and 	XG4980 	(WX8137,WX8762,WX8291);
	and 	XG4981 	(WX8123,WX8762,WX8289);
	and 	XG4982 	(WX8109,WX8762,WX8287);
	and 	XG4983 	(WX8095,WX8762,WX8285);
	and 	XG4984 	(WX8081,WX8762,WX8283);
	and 	XG4985 	(WX8067,WX8762,WX8281);
	and 	XG4986 	(WX8053,WX8762,WX8279);
	and 	XG4987 	(WX8039,WX8762,WX8277);
	and 	XG4988 	(WX8025,WX8762,WX8275);
	and 	XG4989 	(WX8011,WX8762,WX8273);
	and 	XG4990 	(WX7997,WX8762,WX8271);
	and 	XG4991 	(WX7983,WX8762,WX8269);
	and 	XG4992 	(WX7969,WX8762,WX8267);
	and 	XG4993 	(WX7955,WX8762,WX8265);
	and 	XG4994 	(WX7941,WX8762,WX8263);
	and 	XG4995 	(WX7927,WX8762,WX8261);
	and 	XG4996 	(WX7913,WX8762,WX8259);
	and 	XG4997 	(WX7899,WX8762,WX8257);
	and 	XG4998 	(WX7885,WX8762,WX8255);
	and 	XG4999 	(WX7871,WX8762,WX8253);
	and 	XG5000 	(WX7857,WX8762,WX8251);
	and 	XG5001 	(WX7843,WX8762,WX8249);
	and 	XG5002 	(WX7829,WX8762,WX8247);
	and 	XG5003 	(WX7815,WX8762,WX8245);
	and 	XG5004 	(WX7801,WX8762,WX8243);
	nand 	XG5005 	(II22991,II22989,WX7364);
	nand 	XG5006 	(II22960,II22958,WX7362);
	nand 	XG5007 	(II22929,II22927,WX7360);
	nand 	XG5008 	(II22898,II22896,WX7358);
	nand 	XG5009 	(II22867,II22865,WX7356);
	nand 	XG5010 	(II22836,II22834,WX7354);
	nand 	XG5011 	(II22805,II22803,WX7352);
	nand 	XG5012 	(II22774,II22772,WX7350);
	nand 	XG5013 	(II22743,II22741,WX7348);
	nand 	XG5014 	(II22712,II22710,WX7346);
	nand 	XG5015 	(II22681,II22679,WX7344);
	nand 	XG5016 	(II22650,II22648,WX7342);
	nand 	XG5017 	(II22619,II22617,WX7340);
	nand 	XG5018 	(II22588,II22586,WX7338);
	nand 	XG5019 	(II22557,II22555,WX7336);
	nand 	XG5020 	(II22526,II22524,WX7334);
	nand 	XG5021 	(II22495,II22493,WX7332);
	nand 	XG5022 	(II22464,II22462,WX7330);
	nand 	XG5023 	(II22433,II22431,WX7328);
	nand 	XG5024 	(II22402,II22400,WX7326);
	nand 	XG5025 	(II22371,II22369,WX7324);
	nand 	XG5026 	(II22340,II22338,WX7322);
	nand 	XG5027 	(II22309,II22307,WX7320);
	nand 	XG5028 	(II22278,II22276,WX7318);
	nand 	XG5029 	(II22247,II22245,WX7316);
	nand 	XG5030 	(II22216,II22214,WX7314);
	nand 	XG5031 	(II22185,II22183,WX7312);
	nand 	XG5032 	(II22154,II22152,WX7310);
	nand 	XG5033 	(II22123,II22121,WX7308);
	nand 	XG5034 	(II22092,II22090,WX7306);
	nand 	XG5035 	(II22061,II22059,WX7304);
	nand 	XG5036 	(II22030,II22028,WX7302);
	nand 	XG5037 	(II22974,WX7172,WX7467);
	nand 	XG5038 	(II22943,WX7170,WX7467);
	nand 	XG5039 	(II22912,WX7168,WX7467);
	nand 	XG5040 	(II22881,WX7166,WX7467);
	nand 	XG5041 	(II22850,WX7164,WX7467);
	nand 	XG5042 	(II22819,WX7162,WX7467);
	nand 	XG5043 	(II22788,WX7160,WX7467);
	nand 	XG5044 	(II22757,WX7158,WX7467);
	nand 	XG5045 	(II22726,WX7156,WX7467);
	nand 	XG5046 	(II22695,WX7154,WX7467);
	nand 	XG5047 	(II22664,WX7152,WX7467);
	nand 	XG5048 	(II22633,WX7150,WX7467);
	nand 	XG5049 	(II22602,WX7148,WX7467);
	nand 	XG5050 	(II22571,WX7146,WX7467);
	nand 	XG5051 	(II22540,WX7144,WX7467);
	nand 	XG5052 	(II22509,WX7142,WX7467);
	nand 	XG5053 	(II22478,WX7140,WX7466);
	nand 	XG5054 	(II22447,WX7138,WX7466);
	nand 	XG5055 	(II22416,WX7136,WX7466);
	nand 	XG5056 	(II22385,WX7134,WX7466);
	nand 	XG5057 	(II22354,WX7132,WX7466);
	nand 	XG5058 	(II22323,WX7130,WX7466);
	nand 	XG5059 	(II22292,WX7128,WX7466);
	nand 	XG5060 	(II22261,WX7126,WX7466);
	nand 	XG5061 	(II22230,WX7124,WX7466);
	nand 	XG5062 	(II22199,WX7122,WX7466);
	nand 	XG5063 	(II22168,WX7120,WX7466);
	nand 	XG5064 	(II22137,WX7118,WX7466);
	nand 	XG5065 	(II22106,WX7116,WX7466);
	nand 	XG5066 	(II22075,WX7114,WX7466);
	nand 	XG5067 	(II22044,WX7112,WX7466);
	nand 	XG5068 	(II22013,WX7110,WX7466);
	and 	XG5069 	(WX6942,WX7469,WX7012);
	and 	XG5070 	(WX6928,WX7469,WX7010);
	and 	XG5071 	(WX6914,WX7469,WX7008);
	and 	XG5072 	(WX6900,WX7469,WX7006);
	and 	XG5073 	(WX6886,WX7469,WX7004);
	and 	XG5074 	(WX6872,WX7469,WX7002);
	and 	XG5075 	(WX6858,WX7469,WX7000);
	and 	XG5076 	(WX6844,WX7469,WX6998);
	and 	XG5077 	(WX6830,WX7469,WX6996);
	and 	XG5078 	(WX6816,WX7469,WX6994);
	and 	XG5079 	(WX6802,WX7469,WX6992);
	and 	XG5080 	(WX6788,WX7469,WX6990);
	and 	XG5081 	(WX6774,WX7469,WX6988);
	and 	XG5082 	(WX6760,WX7469,WX6986);
	and 	XG5083 	(WX6746,WX7469,WX6984);
	and 	XG5084 	(WX6732,WX7469,WX6982);
	and 	XG5085 	(WX6718,WX7469,WX6980);
	and 	XG5086 	(WX6704,WX7469,WX6978);
	and 	XG5087 	(WX6690,WX7469,WX6976);
	and 	XG5088 	(WX6676,WX7469,WX6974);
	and 	XG5089 	(WX6662,WX7469,WX6972);
	and 	XG5090 	(WX6648,WX7469,WX6970);
	and 	XG5091 	(WX6634,WX7469,WX6968);
	and 	XG5092 	(WX6620,WX7469,WX6966);
	and 	XG5093 	(WX6606,WX7469,WX6964);
	and 	XG5094 	(WX6592,WX7469,WX6962);
	and 	XG5095 	(WX6578,WX7469,WX6960);
	and 	XG5096 	(WX6564,WX7469,WX6958);
	and 	XG5097 	(WX6550,WX7469,WX6956);
	and 	XG5098 	(WX6536,WX7469,WX6954);
	and 	XG5099 	(WX6522,WX7469,WX6952);
	and 	XG5100 	(WX6508,WX7469,WX6950);
	nand 	XG5101 	(II18986,II18984,WX6071);
	nand 	XG5102 	(II18955,II18953,WX6069);
	nand 	XG5103 	(II18924,II18922,WX6067);
	nand 	XG5104 	(II18893,II18891,WX6065);
	nand 	XG5105 	(II18862,II18860,WX6063);
	nand 	XG5106 	(II18831,II18829,WX6061);
	nand 	XG5107 	(II18800,II18798,WX6059);
	nand 	XG5108 	(II18769,II18767,WX6057);
	nand 	XG5109 	(II18738,II18736,WX6055);
	nand 	XG5110 	(II18707,II18705,WX6053);
	nand 	XG5111 	(II18676,II18674,WX6051);
	nand 	XG5112 	(II18645,II18643,WX6049);
	nand 	XG5113 	(II18614,II18612,WX6047);
	nand 	XG5114 	(II18583,II18581,WX6045);
	nand 	XG5115 	(II18552,II18550,WX6043);
	nand 	XG5116 	(II18521,II18519,WX6041);
	nand 	XG5117 	(II18490,II18488,WX6039);
	nand 	XG5118 	(II18459,II18457,WX6037);
	nand 	XG5119 	(II18428,II18426,WX6035);
	nand 	XG5120 	(II18397,II18395,WX6033);
	nand 	XG5121 	(II18366,II18364,WX6031);
	nand 	XG5122 	(II18335,II18333,WX6029);
	nand 	XG5123 	(II18304,II18302,WX6027);
	nand 	XG5124 	(II18273,II18271,WX6025);
	nand 	XG5125 	(II18242,II18240,WX6023);
	nand 	XG5126 	(II18211,II18209,WX6021);
	nand 	XG5127 	(II18180,II18178,WX6019);
	nand 	XG5128 	(II18149,II18147,WX6017);
	nand 	XG5129 	(II18118,II18116,WX6015);
	nand 	XG5130 	(II18087,II18085,WX6013);
	nand 	XG5131 	(II18056,II18054,WX6011);
	nand 	XG5132 	(II18025,II18023,WX6009);
	nand 	XG5133 	(II18969,WX5879,WX6174);
	nand 	XG5134 	(II18938,WX5877,WX6174);
	nand 	XG5135 	(II18907,WX5875,WX6174);
	nand 	XG5136 	(II18876,WX5873,WX6174);
	nand 	XG5137 	(II18845,WX5871,WX6174);
	nand 	XG5138 	(II18814,WX5869,WX6174);
	nand 	XG5139 	(II18783,WX5867,WX6174);
	nand 	XG5140 	(II18752,WX5865,WX6174);
	nand 	XG5141 	(II18721,WX5863,WX6174);
	nand 	XG5142 	(II18690,WX5861,WX6174);
	nand 	XG5143 	(II18659,WX5859,WX6174);
	nand 	XG5144 	(II18628,WX5857,WX6174);
	nand 	XG5145 	(II18597,WX5855,WX6174);
	nand 	XG5146 	(II18566,WX5853,WX6174);
	nand 	XG5147 	(II18535,WX5851,WX6174);
	nand 	XG5148 	(II18504,WX5849,WX6174);
	nand 	XG5149 	(II18473,WX5847,WX6173);
	nand 	XG5150 	(II18442,WX5845,WX6173);
	nand 	XG5151 	(II18411,WX5843,WX6173);
	nand 	XG5152 	(II18380,WX5841,WX6173);
	nand 	XG5153 	(II18349,WX5839,WX6173);
	nand 	XG5154 	(II18318,WX5837,WX6173);
	nand 	XG5155 	(II18287,WX5835,WX6173);
	nand 	XG5156 	(II18256,WX5833,WX6173);
	nand 	XG5157 	(II18225,WX5831,WX6173);
	nand 	XG5158 	(II18194,WX5829,WX6173);
	nand 	XG5159 	(II18163,WX5827,WX6173);
	nand 	XG5160 	(II18132,WX5825,WX6173);
	nand 	XG5161 	(II18101,WX5823,WX6173);
	nand 	XG5162 	(II18070,WX5821,WX6173);
	nand 	XG5163 	(II18039,WX5819,WX6173);
	nand 	XG5164 	(II18008,WX5817,WX6173);
	and 	XG5165 	(WX5649,WX6176,WX5719);
	and 	XG5166 	(WX5635,WX6176,WX5717);
	and 	XG5167 	(WX5621,WX6176,WX5715);
	and 	XG5168 	(WX5607,WX6176,WX5713);
	and 	XG5169 	(WX5593,WX6176,WX5711);
	and 	XG5170 	(WX5579,WX6176,WX5709);
	and 	XG5171 	(WX5565,WX6176,WX5707);
	and 	XG5172 	(WX5551,WX6176,WX5705);
	and 	XG5173 	(WX5537,WX6176,WX5703);
	and 	XG5174 	(WX5523,WX6176,WX5701);
	and 	XG5175 	(WX5509,WX6176,WX5699);
	and 	XG5176 	(WX5495,WX6176,WX5697);
	and 	XG5177 	(WX5481,WX6176,WX5695);
	and 	XG5178 	(WX5467,WX6176,WX5693);
	and 	XG5179 	(WX5453,WX6176,WX5691);
	and 	XG5180 	(WX5439,WX6176,WX5689);
	and 	XG5181 	(WX5425,WX6176,WX5687);
	and 	XG5182 	(WX5411,WX6176,WX5685);
	and 	XG5183 	(WX5397,WX6176,WX5683);
	and 	XG5184 	(WX5383,WX6176,WX5681);
	and 	XG5185 	(WX5369,WX6176,WX5679);
	and 	XG5186 	(WX5355,WX6176,WX5677);
	and 	XG5187 	(WX5341,WX6176,WX5675);
	and 	XG5188 	(WX5327,WX6176,WX5673);
	and 	XG5189 	(WX5313,WX6176,WX5671);
	and 	XG5190 	(WX5299,WX6176,WX5669);
	and 	XG5191 	(WX5285,WX6176,WX5667);
	and 	XG5192 	(WX5271,WX6176,WX5665);
	and 	XG5193 	(WX5257,WX6176,WX5663);
	and 	XG5194 	(WX5243,WX6176,WX5661);
	and 	XG5195 	(WX5229,WX6176,WX5659);
	and 	XG5196 	(WX5215,WX6176,WX5657);
	nand 	XG5197 	(II14981,II14979,WX4778);
	nand 	XG5198 	(II14950,II14948,WX4776);
	nand 	XG5199 	(II14919,II14917,WX4774);
	nand 	XG5200 	(II14888,II14886,WX4772);
	nand 	XG5201 	(II14857,II14855,WX4770);
	nand 	XG5202 	(II14826,II14824,WX4768);
	nand 	XG5203 	(II14795,II14793,WX4766);
	nand 	XG5204 	(II14764,II14762,WX4764);
	nand 	XG5205 	(II14733,II14731,WX4762);
	nand 	XG5206 	(II14702,II14700,WX4760);
	nand 	XG5207 	(II14671,II14669,WX4758);
	nand 	XG5208 	(II14640,II14638,WX4756);
	nand 	XG5209 	(II14609,II14607,WX4754);
	nand 	XG5210 	(II14578,II14576,WX4752);
	nand 	XG5211 	(II14547,II14545,WX4750);
	nand 	XG5212 	(II14516,II14514,WX4748);
	nand 	XG5213 	(II14485,II14483,WX4746);
	nand 	XG5214 	(II14454,II14452,WX4744);
	nand 	XG5215 	(II14423,II14421,WX4742);
	nand 	XG5216 	(II14392,II14390,WX4740);
	nand 	XG5217 	(II14361,II14359,WX4738);
	nand 	XG5218 	(II14330,II14328,WX4736);
	nand 	XG5219 	(II14299,II14297,WX4734);
	nand 	XG5220 	(II14268,II14266,WX4732);
	nand 	XG5221 	(II14237,II14235,WX4730);
	nand 	XG5222 	(II14206,II14204,WX4728);
	nand 	XG5223 	(II14175,II14173,WX4726);
	nand 	XG5224 	(II14144,II14142,WX4724);
	nand 	XG5225 	(II14113,II14111,WX4722);
	nand 	XG5226 	(II14082,II14080,WX4720);
	nand 	XG5227 	(II14051,II14049,WX4718);
	nand 	XG5228 	(II14020,II14018,WX4716);
	nand 	XG5229 	(II14964,WX4586,WX4881);
	nand 	XG5230 	(II14933,WX4584,WX4881);
	nand 	XG5231 	(II14902,WX4582,WX4881);
	nand 	XG5232 	(II14871,WX4580,WX4881);
	nand 	XG5233 	(II14840,WX4578,WX4881);
	nand 	XG5234 	(II14809,WX4576,WX4881);
	nand 	XG5235 	(II14778,WX4574,WX4881);
	nand 	XG5236 	(II14747,WX4572,WX4881);
	nand 	XG5237 	(II14716,WX4570,WX4881);
	nand 	XG5238 	(II14685,WX4568,WX4881);
	nand 	XG5239 	(II14654,WX4566,WX4881);
	nand 	XG5240 	(II14623,WX4564,WX4881);
	nand 	XG5241 	(II14592,WX4562,WX4881);
	nand 	XG5242 	(II14561,WX4560,WX4881);
	nand 	XG5243 	(II14530,WX4558,WX4881);
	nand 	XG5244 	(II14499,WX4556,WX4881);
	nand 	XG5245 	(II14468,WX4554,WX4880);
	nand 	XG5246 	(II14437,WX4552,WX4880);
	nand 	XG5247 	(II14406,WX4550,WX4880);
	nand 	XG5248 	(II14375,WX4548,WX4880);
	nand 	XG5249 	(II14344,WX4546,WX4880);
	nand 	XG5250 	(II14313,WX4544,WX4880);
	nand 	XG5251 	(II14282,WX4542,WX4880);
	nand 	XG5252 	(II14251,WX4540,WX4880);
	nand 	XG5253 	(II14220,WX4538,WX4880);
	nand 	XG5254 	(II14189,WX4536,WX4880);
	nand 	XG5255 	(II14158,WX4534,WX4880);
	nand 	XG5256 	(II14127,WX4532,WX4880);
	nand 	XG5257 	(II14096,WX4530,WX4880);
	nand 	XG5258 	(II14065,WX4528,WX4880);
	nand 	XG5259 	(II14034,WX4526,WX4880);
	nand 	XG5260 	(II14003,WX4524,WX4880);
	and 	XG5261 	(WX4356,WX4883,WX4426);
	and 	XG5262 	(WX4342,WX4883,WX4424);
	and 	XG5263 	(WX4328,WX4883,WX4422);
	and 	XG5264 	(WX4314,WX4883,WX4420);
	and 	XG5265 	(WX4300,WX4883,WX4418);
	and 	XG5266 	(WX4286,WX4883,WX4416);
	and 	XG5267 	(WX4272,WX4883,WX4414);
	and 	XG5268 	(WX4258,WX4883,WX4412);
	and 	XG5269 	(WX4244,WX4883,WX4410);
	and 	XG5270 	(WX4230,WX4883,WX4408);
	and 	XG5271 	(WX4216,WX4883,WX4406);
	and 	XG5272 	(WX4202,WX4883,WX4404);
	and 	XG5273 	(WX4188,WX4883,WX4402);
	and 	XG5274 	(WX4174,WX4883,WX4400);
	and 	XG5275 	(WX4160,WX4883,WX4398);
	and 	XG5276 	(WX4146,WX4883,WX4396);
	and 	XG5277 	(WX4132,WX4883,WX4394);
	and 	XG5278 	(WX4118,WX4883,WX4392);
	and 	XG5279 	(WX4104,WX4883,WX4390);
	and 	XG5280 	(WX4090,WX4883,WX4388);
	and 	XG5281 	(WX4076,WX4883,WX4386);
	and 	XG5282 	(WX4062,WX4883,WX4384);
	and 	XG5283 	(WX4048,WX4883,WX4382);
	and 	XG5284 	(WX4034,WX4883,WX4380);
	and 	XG5285 	(WX4020,WX4883,WX4378);
	and 	XG5286 	(WX4006,WX4883,WX4376);
	and 	XG5287 	(WX3992,WX4883,WX4374);
	and 	XG5288 	(WX3978,WX4883,WX4372);
	and 	XG5289 	(WX3964,WX4883,WX4370);
	and 	XG5290 	(WX3950,WX4883,WX4368);
	and 	XG5291 	(WX3936,WX4883,WX4366);
	and 	XG5292 	(WX3922,WX4883,WX4364);
	nand 	XG5293 	(II10976,II10974,WX3485);
	nand 	XG5294 	(II10945,II10943,WX3483);
	nand 	XG5295 	(II10914,II10912,WX3481);
	nand 	XG5296 	(II10883,II10881,WX3479);
	nand 	XG5297 	(II10852,II10850,WX3477);
	nand 	XG5298 	(II10821,II10819,WX3475);
	nand 	XG5299 	(II10790,II10788,WX3473);
	nand 	XG5300 	(II10759,II10757,WX3471);
	nand 	XG5301 	(II10728,II10726,WX3469);
	nand 	XG5302 	(II10697,II10695,WX3467);
	nand 	XG5303 	(II10666,II10664,WX3465);
	nand 	XG5304 	(II10635,II10633,WX3463);
	nand 	XG5305 	(II10604,II10602,WX3461);
	nand 	XG5306 	(II10573,II10571,WX3459);
	nand 	XG5307 	(II10542,II10540,WX3457);
	nand 	XG5308 	(II10511,II10509,WX3455);
	nand 	XG5309 	(II10480,II10478,WX3453);
	nand 	XG5310 	(II10449,II10447,WX3451);
	nand 	XG5311 	(II10418,II10416,WX3449);
	nand 	XG5312 	(II10387,II10385,WX3447);
	nand 	XG5313 	(II10356,II10354,WX3445);
	nand 	XG5314 	(II10325,II10323,WX3443);
	nand 	XG5315 	(II10294,II10292,WX3441);
	nand 	XG5316 	(II10263,II10261,WX3439);
	nand 	XG5317 	(II10232,II10230,WX3437);
	nand 	XG5318 	(II10201,II10199,WX3435);
	nand 	XG5319 	(II10170,II10168,WX3433);
	nand 	XG5320 	(II10139,II10137,WX3431);
	nand 	XG5321 	(II10108,II10106,WX3429);
	nand 	XG5322 	(II10077,II10075,WX3427);
	nand 	XG5323 	(II10046,II10044,WX3425);
	nand 	XG5324 	(II10015,II10013,WX3423);
	nand 	XG5325 	(II10959,WX3293,WX3588);
	nand 	XG5326 	(II10928,WX3291,WX3588);
	nand 	XG5327 	(II10897,WX3289,WX3588);
	nand 	XG5328 	(II10866,WX3287,WX3588);
	nand 	XG5329 	(II10835,WX3285,WX3588);
	nand 	XG5330 	(II10804,WX3283,WX3588);
	nand 	XG5331 	(II10773,WX3281,WX3588);
	nand 	XG5332 	(II10742,WX3279,WX3588);
	nand 	XG5333 	(II10711,WX3277,WX3588);
	nand 	XG5334 	(II10680,WX3275,WX3588);
	nand 	XG5335 	(II10649,WX3273,WX3588);
	nand 	XG5336 	(II10618,WX3271,WX3588);
	nand 	XG5337 	(II10587,WX3269,WX3588);
	nand 	XG5338 	(II10556,WX3267,WX3588);
	nand 	XG5339 	(II10525,WX3265,WX3588);
	nand 	XG5340 	(II10494,WX3263,WX3588);
	nand 	XG5341 	(II10463,WX3261,WX3587);
	nand 	XG5342 	(II10432,WX3259,WX3587);
	nand 	XG5343 	(II10401,WX3257,WX3587);
	nand 	XG5344 	(II10370,WX3255,WX3587);
	nand 	XG5345 	(II10339,WX3253,WX3587);
	nand 	XG5346 	(II10308,WX3251,WX3587);
	nand 	XG5347 	(II10277,WX3249,WX3587);
	nand 	XG5348 	(II10246,WX3247,WX3587);
	nand 	XG5349 	(II10215,WX3245,WX3587);
	nand 	XG5350 	(II10184,WX3243,WX3587);
	nand 	XG5351 	(II10153,WX3241,WX3587);
	nand 	XG5352 	(II10122,WX3239,WX3587);
	nand 	XG5353 	(II10091,WX3237,WX3587);
	nand 	XG5354 	(II10060,WX3235,WX3587);
	nand 	XG5355 	(II10029,WX3233,WX3587);
	nand 	XG5356 	(II9998,WX3231,WX3587);
	and 	XG5357 	(WX3063,WX3590,WX3133);
	and 	XG5358 	(WX3049,WX3590,WX3131);
	and 	XG5359 	(WX3035,WX3590,WX3129);
	and 	XG5360 	(WX3021,WX3590,WX3127);
	and 	XG5361 	(WX3007,WX3590,WX3125);
	and 	XG5362 	(WX2993,WX3590,WX3123);
	and 	XG5363 	(WX2979,WX3590,WX3121);
	and 	XG5364 	(WX2965,WX3590,WX3119);
	and 	XG5365 	(WX2951,WX3590,WX3117);
	and 	XG5366 	(WX2937,WX3590,WX3115);
	and 	XG5367 	(WX2923,WX3590,WX3113);
	and 	XG5368 	(WX2909,WX3590,WX3111);
	and 	XG5369 	(WX2895,WX3590,WX3109);
	and 	XG5370 	(WX2881,WX3590,WX3107);
	and 	XG5371 	(WX2867,WX3590,WX3105);
	and 	XG5372 	(WX2853,WX3590,WX3103);
	and 	XG5373 	(WX2839,WX3590,WX3101);
	and 	XG5374 	(WX2825,WX3590,WX3099);
	and 	XG5375 	(WX2811,WX3590,WX3097);
	and 	XG5376 	(WX2797,WX3590,WX3095);
	and 	XG5377 	(WX2783,WX3590,WX3093);
	and 	XG5378 	(WX2769,WX3590,WX3091);
	and 	XG5379 	(WX2755,WX3590,WX3089);
	and 	XG5380 	(WX2741,WX3590,WX3087);
	and 	XG5381 	(WX2727,WX3590,WX3085);
	and 	XG5382 	(WX2713,WX3590,WX3083);
	and 	XG5383 	(WX2699,WX3590,WX3081);
	and 	XG5384 	(WX2685,WX3590,WX3079);
	and 	XG5385 	(WX2671,WX3590,WX3077);
	and 	XG5386 	(WX2657,WX3590,WX3075);
	and 	XG5387 	(WX2643,WX3590,WX3073);
	and 	XG5388 	(WX2629,WX3590,WX3071);
	nand 	XG5389 	(II6971,II6969,WX2192);
	nand 	XG5390 	(II6940,II6938,WX2190);
	nand 	XG5391 	(II6909,II6907,WX2188);
	nand 	XG5392 	(II6878,II6876,WX2186);
	nand 	XG5393 	(II6847,II6845,WX2184);
	nand 	XG5394 	(II6816,II6814,WX2182);
	nand 	XG5395 	(II6785,II6783,WX2180);
	nand 	XG5396 	(II6754,II6752,WX2178);
	nand 	XG5397 	(II6723,II6721,WX2176);
	nand 	XG5398 	(II6692,II6690,WX2174);
	nand 	XG5399 	(II6661,II6659,WX2172);
	nand 	XG5400 	(II6630,II6628,WX2170);
	nand 	XG5401 	(II6599,II6597,WX2168);
	nand 	XG5402 	(II6568,II6566,WX2166);
	nand 	XG5403 	(II6537,II6535,WX2164);
	nand 	XG5404 	(II6506,II6504,WX2162);
	nand 	XG5405 	(II6475,II6473,WX2160);
	nand 	XG5406 	(II6444,II6442,WX2158);
	nand 	XG5407 	(II6413,II6411,WX2156);
	nand 	XG5408 	(II6382,II6380,WX2154);
	nand 	XG5409 	(II6351,II6349,WX2152);
	nand 	XG5410 	(II6320,II6318,WX2150);
	nand 	XG5411 	(II6289,II6287,WX2148);
	nand 	XG5412 	(II6258,II6256,WX2146);
	nand 	XG5413 	(II6227,II6225,WX2144);
	nand 	XG5414 	(II6196,II6194,WX2142);
	nand 	XG5415 	(II6165,II6163,WX2140);
	nand 	XG5416 	(II6134,II6132,WX2138);
	nand 	XG5417 	(II6103,II6101,WX2136);
	nand 	XG5418 	(II6072,II6070,WX2134);
	nand 	XG5419 	(II6041,II6039,WX2132);
	nand 	XG5420 	(II6010,II6008,WX2130);
	nand 	XG5421 	(II6954,WX2000,WX2295);
	nand 	XG5422 	(II6923,WX1998,WX2295);
	nand 	XG5423 	(II6892,WX1996,WX2295);
	nand 	XG5424 	(II6861,WX1994,WX2295);
	nand 	XG5425 	(II6830,WX1992,WX2295);
	nand 	XG5426 	(II6799,WX1990,WX2295);
	nand 	XG5427 	(II6768,WX1988,WX2295);
	nand 	XG5428 	(II6737,WX1986,WX2295);
	nand 	XG5429 	(II6706,WX1984,WX2295);
	nand 	XG5430 	(II6675,WX1982,WX2295);
	nand 	XG5431 	(II6644,WX1980,WX2295);
	nand 	XG5432 	(II6613,WX1978,WX2295);
	nand 	XG5433 	(II6582,WX1976,WX2295);
	nand 	XG5434 	(II6551,WX1974,WX2295);
	nand 	XG5435 	(II6520,WX1972,WX2295);
	nand 	XG5436 	(II6489,WX1970,WX2295);
	nand 	XG5437 	(II6458,WX1968,WX2294);
	nand 	XG5438 	(II6427,WX1966,WX2294);
	nand 	XG5439 	(II6396,WX1964,WX2294);
	nand 	XG5440 	(II6365,WX1962,WX2294);
	nand 	XG5441 	(II6334,WX1960,WX2294);
	nand 	XG5442 	(II6303,WX1958,WX2294);
	nand 	XG5443 	(II6272,WX1956,WX2294);
	nand 	XG5444 	(II6241,WX1954,WX2294);
	nand 	XG5445 	(II6210,WX1952,WX2294);
	nand 	XG5446 	(II6179,WX1950,WX2294);
	nand 	XG5447 	(II6148,WX1948,WX2294);
	nand 	XG5448 	(II6117,WX1946,WX2294);
	nand 	XG5449 	(II6086,WX1944,WX2294);
	nand 	XG5450 	(II6055,WX1942,WX2294);
	nand 	XG5451 	(II6024,WX1940,WX2294);
	nand 	XG5452 	(II5993,WX1938,WX2294);
	and 	XG5453 	(WX1770,WX2297,WX1840);
	and 	XG5454 	(WX1756,WX2297,WX1838);
	and 	XG5455 	(WX1742,WX2297,WX1836);
	and 	XG5456 	(WX1728,WX2297,WX1834);
	and 	XG5457 	(WX1714,WX2297,WX1832);
	and 	XG5458 	(WX1700,WX2297,WX1830);
	and 	XG5459 	(WX1686,WX2297,WX1828);
	and 	XG5460 	(WX1672,WX2297,WX1826);
	and 	XG5461 	(WX1658,WX2297,WX1824);
	and 	XG5462 	(WX1644,WX2297,WX1822);
	and 	XG5463 	(WX1630,WX2297,WX1820);
	and 	XG5464 	(WX1616,WX2297,WX1818);
	and 	XG5465 	(WX1602,WX2297,WX1816);
	and 	XG5466 	(WX1588,WX2297,WX1814);
	and 	XG5467 	(WX1574,WX2297,WX1812);
	and 	XG5468 	(WX1560,WX2297,WX1810);
	and 	XG5469 	(WX1546,WX2297,WX1808);
	and 	XG5470 	(WX1532,WX2297,WX1806);
	and 	XG5471 	(WX1518,WX2297,WX1804);
	and 	XG5472 	(WX1504,WX2297,WX1802);
	and 	XG5473 	(WX1490,WX2297,WX1800);
	and 	XG5474 	(WX1476,WX2297,WX1798);
	and 	XG5475 	(WX1462,WX2297,WX1796);
	and 	XG5476 	(WX1448,WX2297,WX1794);
	and 	XG5477 	(WX1434,WX2297,WX1792);
	and 	XG5478 	(WX1420,WX2297,WX1790);
	and 	XG5479 	(WX1406,WX2297,WX1788);
	and 	XG5480 	(WX1392,WX2297,WX1786);
	and 	XG5481 	(WX1378,WX2297,WX1784);
	and 	XG5482 	(WX1364,WX2297,WX1782);
	and 	XG5483 	(WX1350,WX2297,WX1780);
	and 	XG5484 	(WX1336,WX2297,WX1778);
	nand 	XG5485 	(II2966,II2964,WX899);
	nand 	XG5486 	(II2935,II2933,WX897);
	nand 	XG5487 	(II2904,II2902,WX895);
	nand 	XG5488 	(II2873,II2871,WX893);
	nand 	XG5489 	(II2842,II2840,WX891);
	nand 	XG5490 	(II2811,II2809,WX889);
	nand 	XG5491 	(II2780,II2778,WX887);
	nand 	XG5492 	(II2749,II2747,WX885);
	nand 	XG5493 	(II2718,II2716,WX883);
	nand 	XG5494 	(II2687,II2685,WX881);
	nand 	XG5495 	(II2656,II2654,WX879);
	nand 	XG5496 	(II2625,II2623,WX877);
	nand 	XG5497 	(II2594,II2592,WX875);
	nand 	XG5498 	(II2563,II2561,WX873);
	nand 	XG5499 	(II2532,II2530,WX871);
	nand 	XG5500 	(II2501,II2499,WX869);
	nand 	XG5501 	(II2470,II2468,WX867);
	nand 	XG5502 	(II2439,II2437,WX865);
	nand 	XG5503 	(II2408,II2406,WX863);
	nand 	XG5504 	(II2377,II2375,WX861);
	nand 	XG5505 	(II2346,II2344,WX859);
	nand 	XG5506 	(II2315,II2313,WX857);
	nand 	XG5507 	(II2284,II2282,WX855);
	nand 	XG5508 	(II2253,II2251,WX853);
	nand 	XG5509 	(II2222,II2220,WX851);
	nand 	XG5510 	(II2191,II2189,WX849);
	nand 	XG5511 	(II2160,II2158,WX847);
	nand 	XG5512 	(II2129,II2127,WX845);
	nand 	XG5513 	(II2098,II2096,WX843);
	nand 	XG5514 	(II2067,II2065,WX841);
	nand 	XG5515 	(II2036,II2034,WX839);
	nand 	XG5516 	(II2005,II2003,WX837);
	nand 	XG5517 	(II2949,WX707,WX1002);
	nand 	XG5518 	(II2918,WX705,WX1002);
	nand 	XG5519 	(II2887,WX703,WX1002);
	nand 	XG5520 	(II2856,WX701,WX1002);
	nand 	XG5521 	(II2825,WX699,WX1002);
	nand 	XG5522 	(II2794,WX697,WX1002);
	nand 	XG5523 	(II2763,WX695,WX1002);
	nand 	XG5524 	(II2732,WX693,WX1002);
	nand 	XG5525 	(II2701,WX691,WX1002);
	nand 	XG5526 	(II2670,WX689,WX1002);
	nand 	XG5527 	(II2639,WX687,WX1002);
	nand 	XG5528 	(II2608,WX685,WX1002);
	nand 	XG5529 	(II2577,WX683,WX1002);
	nand 	XG5530 	(II2546,WX681,WX1002);
	nand 	XG5531 	(II2515,WX679,WX1002);
	nand 	XG5532 	(II2484,WX677,WX1002);
	nand 	XG5533 	(II2453,WX675,WX1001);
	nand 	XG5534 	(II2422,WX673,WX1001);
	nand 	XG5535 	(II2391,WX671,WX1001);
	nand 	XG5536 	(II2360,WX669,WX1001);
	nand 	XG5537 	(II2329,WX667,WX1001);
	nand 	XG5538 	(II2298,WX665,WX1001);
	nand 	XG5539 	(II2267,WX663,WX1001);
	nand 	XG5540 	(II2236,WX661,WX1001);
	nand 	XG5541 	(II2205,WX659,WX1001);
	nand 	XG5542 	(II2174,WX657,WX1001);
	nand 	XG5543 	(II2143,WX655,WX1001);
	nand 	XG5544 	(II2112,WX653,WX1001);
	nand 	XG5545 	(II2081,WX651,WX1001);
	nand 	XG5546 	(II2050,WX649,WX1001);
	nand 	XG5547 	(II2019,WX647,WX1001);
	nand 	XG5548 	(II1988,WX645,WX1001);
	and 	XG5549 	(WX477,WX1004,WX547);
	and 	XG5550 	(WX463,WX1004,WX545);
	and 	XG5551 	(WX449,WX1004,WX543);
	and 	XG5552 	(WX435,WX1004,WX541);
	and 	XG5553 	(WX421,WX1004,WX539);
	and 	XG5554 	(WX407,WX1004,WX537);
	and 	XG5555 	(WX393,WX1004,WX535);
	and 	XG5556 	(WX379,WX1004,WX533);
	and 	XG5557 	(WX365,WX1004,WX531);
	and 	XG5558 	(WX351,WX1004,WX529);
	and 	XG5559 	(WX337,WX1004,WX527);
	and 	XG5560 	(WX323,WX1004,WX525);
	and 	XG5561 	(WX309,WX1004,WX523);
	and 	XG5562 	(WX295,WX1004,WX521);
	and 	XG5563 	(WX281,WX1004,WX519);
	and 	XG5564 	(WX267,WX1004,WX517);
	and 	XG5565 	(WX253,WX1004,WX515);
	and 	XG5566 	(WX239,WX1004,WX513);
	and 	XG5567 	(WX225,WX1004,WX511);
	and 	XG5568 	(WX211,WX1004,WX509);
	and 	XG5569 	(WX197,WX1004,WX507);
	and 	XG5570 	(WX183,WX1004,WX505);
	and 	XG5571 	(WX169,WX1004,WX503);
	and 	XG5572 	(WX155,WX1004,WX501);
	and 	XG5573 	(WX141,WX1004,WX499);
	and 	XG5574 	(WX127,WX1004,WX497);
	and 	XG5575 	(WX113,WX1004,WX495);
	and 	XG5576 	(WX99,WX1004,WX493);
	and 	XG5577 	(WX85,WX1004,WX491);
	and 	XG5578 	(WX71,WX1004,WX489);
	and 	XG5579 	(WX57,WX1004,WX487);
	and 	XG5580 	(WX43,WX1004,WX485);
	and 	XG5581 	(WX10383,WX11348,CRC_OUT_1_31);
	and 	XG5582 	(WX10397,WX11348,CRC_OUT_1_30);
	and 	XG5583 	(WX10411,WX11348,CRC_OUT_1_29);
	and 	XG5584 	(WX10425,WX11348,CRC_OUT_1_28);
	and 	XG5585 	(WX10439,WX11348,CRC_OUT_1_27);
	and 	XG5586 	(WX10453,WX11348,CRC_OUT_1_26);
	and 	XG5587 	(WX10467,WX11348,CRC_OUT_1_25);
	and 	XG5588 	(WX10481,WX11348,CRC_OUT_1_24);
	and 	XG5589 	(WX10495,WX11348,CRC_OUT_1_23);
	and 	XG5590 	(WX10509,WX11348,CRC_OUT_1_22);
	and 	XG5591 	(WX10523,WX11348,CRC_OUT_1_21);
	and 	XG5592 	(WX10537,WX11348,CRC_OUT_1_20);
	and 	XG5593 	(WX10551,WX11348,CRC_OUT_1_19);
	and 	XG5594 	(WX10565,WX11348,CRC_OUT_1_18);
	and 	XG5595 	(WX10579,WX11348,CRC_OUT_1_17);
	and 	XG5596 	(WX10593,WX11348,CRC_OUT_1_16);
	and 	XG5597 	(WX10607,WX11348,CRC_OUT_1_15);
	and 	XG5598 	(WX10621,WX11348,CRC_OUT_1_14);
	and 	XG5599 	(WX10635,WX11348,CRC_OUT_1_13);
	and 	XG5600 	(WX10649,WX11348,CRC_OUT_1_12);
	and 	XG5601 	(WX10663,WX11348,CRC_OUT_1_11);
	and 	XG5602 	(WX10677,WX11348,CRC_OUT_1_10);
	and 	XG5603 	(WX10691,WX11348,CRC_OUT_1_9);
	and 	XG5604 	(WX10705,WX11348,CRC_OUT_1_8);
	and 	XG5605 	(WX10719,WX11348,CRC_OUT_1_7);
	and 	XG5606 	(WX10733,WX11348,CRC_OUT_1_6);
	and 	XG5607 	(WX10747,WX11348,CRC_OUT_1_5);
	and 	XG5608 	(WX10761,WX11348,CRC_OUT_1_4);
	and 	XG5609 	(WX10775,WX11348,CRC_OUT_1_3);
	and 	XG5610 	(WX10789,WX11348,CRC_OUT_1_2);
	and 	XG5611 	(WX10803,WX11348,CRC_OUT_1_1);
	and 	XG5612 	(WX10817,WX11348,CRC_OUT_1_0);
	and 	XG5613 	(WX9090,WX10055,CRC_OUT_2_31);
	and 	XG5614 	(WX9104,WX10055,CRC_OUT_2_30);
	and 	XG5615 	(WX9118,WX10055,CRC_OUT_2_29);
	and 	XG5616 	(WX9132,WX10055,CRC_OUT_2_28);
	and 	XG5617 	(WX9146,WX10055,CRC_OUT_2_27);
	and 	XG5618 	(WX9160,WX10055,CRC_OUT_2_26);
	and 	XG5619 	(WX9174,WX10055,CRC_OUT_2_25);
	and 	XG5620 	(WX9188,WX10055,CRC_OUT_2_24);
	and 	XG5621 	(WX9202,WX10055,CRC_OUT_2_23);
	and 	XG5622 	(WX9216,WX10055,CRC_OUT_2_22);
	and 	XG5623 	(WX9230,WX10055,CRC_OUT_2_21);
	and 	XG5624 	(WX9244,WX10055,CRC_OUT_2_20);
	and 	XG5625 	(WX9258,WX10055,CRC_OUT_2_19);
	and 	XG5626 	(WX9272,WX10055,CRC_OUT_2_18);
	and 	XG5627 	(WX9286,WX10055,CRC_OUT_2_17);
	and 	XG5628 	(WX9300,WX10055,CRC_OUT_2_16);
	and 	XG5629 	(WX9314,WX10055,CRC_OUT_2_15);
	and 	XG5630 	(WX9328,WX10055,CRC_OUT_2_14);
	and 	XG5631 	(WX9342,WX10055,CRC_OUT_2_13);
	and 	XG5632 	(WX9356,WX10055,CRC_OUT_2_12);
	and 	XG5633 	(WX9370,WX10055,CRC_OUT_2_11);
	and 	XG5634 	(WX9384,WX10055,CRC_OUT_2_10);
	and 	XG5635 	(WX9398,WX10055,CRC_OUT_2_9);
	and 	XG5636 	(WX9412,WX10055,CRC_OUT_2_8);
	and 	XG5637 	(WX9426,WX10055,CRC_OUT_2_7);
	and 	XG5638 	(WX9440,WX10055,CRC_OUT_2_6);
	and 	XG5639 	(WX9454,WX10055,CRC_OUT_2_5);
	and 	XG5640 	(WX9468,WX10055,CRC_OUT_2_4);
	and 	XG5641 	(WX9482,WX10055,CRC_OUT_2_3);
	and 	XG5642 	(WX9496,WX10055,CRC_OUT_2_2);
	and 	XG5643 	(WX9510,WX10055,CRC_OUT_2_1);
	and 	XG5644 	(WX9524,WX10055,CRC_OUT_2_0);
	and 	XG5645 	(WX7797,WX8762,CRC_OUT_3_31);
	and 	XG5646 	(WX7811,WX8762,CRC_OUT_3_30);
	and 	XG5647 	(WX7825,WX8762,CRC_OUT_3_29);
	and 	XG5648 	(WX7839,WX8762,CRC_OUT_3_28);
	and 	XG5649 	(WX7853,WX8762,CRC_OUT_3_27);
	and 	XG5650 	(WX7867,WX8762,CRC_OUT_3_26);
	and 	XG5651 	(WX7881,WX8762,CRC_OUT_3_25);
	and 	XG5652 	(WX7895,WX8762,CRC_OUT_3_24);
	and 	XG5653 	(WX7909,WX8762,CRC_OUT_3_23);
	and 	XG5654 	(WX7923,WX8762,CRC_OUT_3_22);
	and 	XG5655 	(WX7937,WX8762,CRC_OUT_3_21);
	and 	XG5656 	(WX7951,WX8762,CRC_OUT_3_20);
	and 	XG5657 	(WX7965,WX8762,CRC_OUT_3_19);
	and 	XG5658 	(WX7979,WX8762,CRC_OUT_3_18);
	and 	XG5659 	(WX7993,WX8762,CRC_OUT_3_17);
	and 	XG5660 	(WX8007,WX8762,CRC_OUT_3_16);
	and 	XG5661 	(WX8021,WX8762,CRC_OUT_3_15);
	and 	XG5662 	(WX8035,WX8762,CRC_OUT_3_14);
	and 	XG5663 	(WX8049,WX8762,CRC_OUT_3_13);
	and 	XG5664 	(WX8063,WX8762,CRC_OUT_3_12);
	and 	XG5665 	(WX8077,WX8762,CRC_OUT_3_11);
	and 	XG5666 	(WX8091,WX8762,CRC_OUT_3_10);
	and 	XG5667 	(WX8105,WX8762,CRC_OUT_3_9);
	and 	XG5668 	(WX8119,WX8762,CRC_OUT_3_8);
	and 	XG5669 	(WX8133,WX8762,CRC_OUT_3_7);
	and 	XG5670 	(WX8147,WX8762,CRC_OUT_3_6);
	and 	XG5671 	(WX8161,WX8762,CRC_OUT_3_5);
	and 	XG5672 	(WX8175,WX8762,CRC_OUT_3_4);
	and 	XG5673 	(WX8189,WX8762,CRC_OUT_3_3);
	and 	XG5674 	(WX8203,WX8762,CRC_OUT_3_2);
	and 	XG5675 	(WX8217,WX8762,CRC_OUT_3_1);
	and 	XG5676 	(WX8231,WX8762,CRC_OUT_3_0);
	and 	XG5677 	(WX6504,WX7469,CRC_OUT_4_31);
	and 	XG5678 	(WX6518,WX7469,CRC_OUT_4_30);
	and 	XG5679 	(WX6532,WX7469,CRC_OUT_4_29);
	and 	XG5680 	(WX6546,WX7469,CRC_OUT_4_28);
	and 	XG5681 	(WX6560,WX7469,CRC_OUT_4_27);
	and 	XG5682 	(WX6574,WX7469,CRC_OUT_4_26);
	and 	XG5683 	(WX6588,WX7469,CRC_OUT_4_25);
	and 	XG5684 	(WX6602,WX7469,CRC_OUT_4_24);
	and 	XG5685 	(WX6616,WX7469,CRC_OUT_4_23);
	and 	XG5686 	(WX6630,WX7469,CRC_OUT_4_22);
	and 	XG5687 	(WX6644,WX7469,CRC_OUT_4_21);
	and 	XG5688 	(WX6658,WX7469,CRC_OUT_4_20);
	and 	XG5689 	(WX6672,WX7469,CRC_OUT_4_19);
	and 	XG5690 	(WX6686,WX7469,CRC_OUT_4_18);
	and 	XG5691 	(WX6700,WX7469,CRC_OUT_4_17);
	and 	XG5692 	(WX6714,WX7469,CRC_OUT_4_16);
	and 	XG5693 	(WX6728,WX7469,CRC_OUT_4_15);
	and 	XG5694 	(WX6742,WX7469,CRC_OUT_4_14);
	and 	XG5695 	(WX6756,WX7469,CRC_OUT_4_13);
	and 	XG5696 	(WX6770,WX7469,CRC_OUT_4_12);
	and 	XG5697 	(WX6784,WX7469,CRC_OUT_4_11);
	and 	XG5698 	(WX6798,WX7469,CRC_OUT_4_10);
	and 	XG5699 	(WX6812,WX7469,CRC_OUT_4_9);
	and 	XG5700 	(WX6826,WX7469,CRC_OUT_4_8);
	and 	XG5701 	(WX6840,WX7469,CRC_OUT_4_7);
	and 	XG5702 	(WX6854,WX7469,CRC_OUT_4_6);
	and 	XG5703 	(WX6868,WX7469,CRC_OUT_4_5);
	and 	XG5704 	(WX6882,WX7469,CRC_OUT_4_4);
	and 	XG5705 	(WX6896,WX7469,CRC_OUT_4_3);
	and 	XG5706 	(WX6910,WX7469,CRC_OUT_4_2);
	and 	XG5707 	(WX6924,WX7469,CRC_OUT_4_1);
	and 	XG5708 	(WX6938,WX7469,CRC_OUT_4_0);
	and 	XG5709 	(WX5211,WX6176,CRC_OUT_5_31);
	and 	XG5710 	(WX5225,WX6176,CRC_OUT_5_30);
	and 	XG5711 	(WX5239,WX6176,CRC_OUT_5_29);
	and 	XG5712 	(WX5253,WX6176,CRC_OUT_5_28);
	and 	XG5713 	(WX5267,WX6176,CRC_OUT_5_27);
	and 	XG5714 	(WX5281,WX6176,CRC_OUT_5_26);
	and 	XG5715 	(WX5295,WX6176,CRC_OUT_5_25);
	and 	XG5716 	(WX5309,WX6176,CRC_OUT_5_24);
	and 	XG5717 	(WX5323,WX6176,CRC_OUT_5_23);
	and 	XG5718 	(WX5337,WX6176,CRC_OUT_5_22);
	and 	XG5719 	(WX5351,WX6176,CRC_OUT_5_21);
	and 	XG5720 	(WX5365,WX6176,CRC_OUT_5_20);
	and 	XG5721 	(WX5379,WX6176,CRC_OUT_5_19);
	and 	XG5722 	(WX5393,WX6176,CRC_OUT_5_18);
	and 	XG5723 	(WX5407,WX6176,CRC_OUT_5_17);
	and 	XG5724 	(WX5421,WX6176,CRC_OUT_5_16);
	and 	XG5725 	(WX5435,WX6176,CRC_OUT_5_15);
	and 	XG5726 	(WX5449,WX6176,CRC_OUT_5_14);
	and 	XG5727 	(WX5463,WX6176,CRC_OUT_5_13);
	and 	XG5728 	(WX5477,WX6176,CRC_OUT_5_12);
	and 	XG5729 	(WX5491,WX6176,CRC_OUT_5_11);
	and 	XG5730 	(WX5505,WX6176,CRC_OUT_5_10);
	and 	XG5731 	(WX5519,WX6176,CRC_OUT_5_9);
	and 	XG5732 	(WX5533,WX6176,CRC_OUT_5_8);
	and 	XG5733 	(WX5547,WX6176,CRC_OUT_5_7);
	and 	XG5734 	(WX5561,WX6176,CRC_OUT_5_6);
	and 	XG5735 	(WX5575,WX6176,CRC_OUT_5_5);
	and 	XG5736 	(WX5589,WX6176,CRC_OUT_5_4);
	and 	XG5737 	(WX5603,WX6176,CRC_OUT_5_3);
	and 	XG5738 	(WX5617,WX6176,CRC_OUT_5_2);
	and 	XG5739 	(WX5631,WX6176,CRC_OUT_5_1);
	and 	XG5740 	(WX5645,WX6176,CRC_OUT_5_0);
	and 	XG5741 	(WX3918,WX4883,CRC_OUT_6_31);
	and 	XG5742 	(WX3932,WX4883,CRC_OUT_6_30);
	and 	XG5743 	(WX3946,WX4883,CRC_OUT_6_29);
	and 	XG5744 	(WX3960,WX4883,CRC_OUT_6_28);
	and 	XG5745 	(WX3974,WX4883,CRC_OUT_6_27);
	and 	XG5746 	(WX3988,WX4883,CRC_OUT_6_26);
	and 	XG5747 	(WX4002,WX4883,CRC_OUT_6_25);
	and 	XG5748 	(WX4016,WX4883,CRC_OUT_6_24);
	and 	XG5749 	(WX4030,WX4883,CRC_OUT_6_23);
	and 	XG5750 	(WX4044,WX4883,CRC_OUT_6_22);
	and 	XG5751 	(WX4058,WX4883,CRC_OUT_6_21);
	and 	XG5752 	(WX4072,WX4883,CRC_OUT_6_20);
	and 	XG5753 	(WX4086,WX4883,CRC_OUT_6_19);
	and 	XG5754 	(WX4100,WX4883,CRC_OUT_6_18);
	and 	XG5755 	(WX4114,WX4883,CRC_OUT_6_17);
	and 	XG5756 	(WX4128,WX4883,CRC_OUT_6_16);
	and 	XG5757 	(WX4142,WX4883,CRC_OUT_6_15);
	and 	XG5758 	(WX4156,WX4883,CRC_OUT_6_14);
	and 	XG5759 	(WX4170,WX4883,CRC_OUT_6_13);
	and 	XG5760 	(WX4184,WX4883,CRC_OUT_6_12);
	and 	XG5761 	(WX4198,WX4883,CRC_OUT_6_11);
	and 	XG5762 	(WX4212,WX4883,CRC_OUT_6_10);
	and 	XG5763 	(WX4226,WX4883,CRC_OUT_6_9);
	and 	XG5764 	(WX4240,WX4883,CRC_OUT_6_8);
	and 	XG5765 	(WX4254,WX4883,CRC_OUT_6_7);
	and 	XG5766 	(WX4268,WX4883,CRC_OUT_6_6);
	and 	XG5767 	(WX4282,WX4883,CRC_OUT_6_5);
	and 	XG5768 	(WX4296,WX4883,CRC_OUT_6_4);
	and 	XG5769 	(WX4310,WX4883,CRC_OUT_6_3);
	and 	XG5770 	(WX4324,WX4883,CRC_OUT_6_2);
	and 	XG5771 	(WX4338,WX4883,CRC_OUT_6_1);
	and 	XG5772 	(WX4352,WX4883,CRC_OUT_6_0);
	and 	XG5773 	(WX2625,WX3590,CRC_OUT_7_31);
	and 	XG5774 	(WX2639,WX3590,CRC_OUT_7_30);
	and 	XG5775 	(WX2653,WX3590,CRC_OUT_7_29);
	and 	XG5776 	(WX2667,WX3590,CRC_OUT_7_28);
	and 	XG5777 	(WX2681,WX3590,CRC_OUT_7_27);
	and 	XG5778 	(WX2695,WX3590,CRC_OUT_7_26);
	and 	XG5779 	(WX2709,WX3590,CRC_OUT_7_25);
	and 	XG5780 	(WX2723,WX3590,CRC_OUT_7_24);
	and 	XG5781 	(WX2737,WX3590,CRC_OUT_7_23);
	and 	XG5782 	(WX2751,WX3590,CRC_OUT_7_22);
	and 	XG5783 	(WX2765,WX3590,CRC_OUT_7_21);
	and 	XG5784 	(WX2779,WX3590,CRC_OUT_7_20);
	and 	XG5785 	(WX2793,WX3590,CRC_OUT_7_19);
	and 	XG5786 	(WX2807,WX3590,CRC_OUT_7_18);
	and 	XG5787 	(WX2821,WX3590,CRC_OUT_7_17);
	and 	XG5788 	(WX2835,WX3590,CRC_OUT_7_16);
	and 	XG5789 	(WX2849,WX3590,CRC_OUT_7_15);
	and 	XG5790 	(WX2863,WX3590,CRC_OUT_7_14);
	and 	XG5791 	(WX2877,WX3590,CRC_OUT_7_13);
	and 	XG5792 	(WX2891,WX3590,CRC_OUT_7_12);
	and 	XG5793 	(WX2905,WX3590,CRC_OUT_7_11);
	and 	XG5794 	(WX2919,WX3590,CRC_OUT_7_10);
	and 	XG5795 	(WX2933,WX3590,CRC_OUT_7_9);
	and 	XG5796 	(WX2947,WX3590,CRC_OUT_7_8);
	and 	XG5797 	(WX2961,WX3590,CRC_OUT_7_7);
	and 	XG5798 	(WX2975,WX3590,CRC_OUT_7_6);
	and 	XG5799 	(WX2989,WX3590,CRC_OUT_7_5);
	and 	XG5800 	(WX3003,WX3590,CRC_OUT_7_4);
	and 	XG5801 	(WX3017,WX3590,CRC_OUT_7_3);
	and 	XG5802 	(WX3031,WX3590,CRC_OUT_7_2);
	and 	XG5803 	(WX3045,WX3590,CRC_OUT_7_1);
	and 	XG5804 	(WX3059,WX3590,CRC_OUT_7_0);
	and 	XG5805 	(WX1332,WX2297,CRC_OUT_8_31);
	and 	XG5806 	(WX1346,WX2297,CRC_OUT_8_30);
	and 	XG5807 	(WX1360,WX2297,CRC_OUT_8_29);
	and 	XG5808 	(WX1374,WX2297,CRC_OUT_8_28);
	and 	XG5809 	(WX1388,WX2297,CRC_OUT_8_27);
	and 	XG5810 	(WX1402,WX2297,CRC_OUT_8_26);
	and 	XG5811 	(WX1416,WX2297,CRC_OUT_8_25);
	and 	XG5812 	(WX1430,WX2297,CRC_OUT_8_24);
	and 	XG5813 	(WX1444,WX2297,CRC_OUT_8_23);
	and 	XG5814 	(WX1458,WX2297,CRC_OUT_8_22);
	and 	XG5815 	(WX1472,WX2297,CRC_OUT_8_21);
	and 	XG5816 	(WX1486,WX2297,CRC_OUT_8_20);
	and 	XG5817 	(WX1500,WX2297,CRC_OUT_8_19);
	and 	XG5818 	(WX1514,WX2297,CRC_OUT_8_18);
	and 	XG5819 	(WX1528,WX2297,CRC_OUT_8_17);
	and 	XG5820 	(WX1542,WX2297,CRC_OUT_8_16);
	and 	XG5821 	(WX1556,WX2297,CRC_OUT_8_15);
	and 	XG5822 	(WX1570,WX2297,CRC_OUT_8_14);
	and 	XG5823 	(WX1584,WX2297,CRC_OUT_8_13);
	and 	XG5824 	(WX1598,WX2297,CRC_OUT_8_12);
	and 	XG5825 	(WX1612,WX2297,CRC_OUT_8_11);
	and 	XG5826 	(WX1626,WX2297,CRC_OUT_8_10);
	and 	XG5827 	(WX1640,WX2297,CRC_OUT_8_9);
	and 	XG5828 	(WX1654,WX2297,CRC_OUT_8_8);
	and 	XG5829 	(WX1668,WX2297,CRC_OUT_8_7);
	and 	XG5830 	(WX1682,WX2297,CRC_OUT_8_6);
	and 	XG5831 	(WX1696,WX2297,CRC_OUT_8_5);
	and 	XG5832 	(WX1710,WX2297,CRC_OUT_8_4);
	and 	XG5833 	(WX1724,WX2297,CRC_OUT_8_3);
	and 	XG5834 	(WX1738,WX2297,CRC_OUT_8_2);
	and 	XG5835 	(WX1752,WX2297,CRC_OUT_8_1);
	and 	XG5836 	(WX1766,WX2297,CRC_OUT_8_0);
	and 	XG5837 	(WX39,WX1004,CRC_OUT_9_31);
	and 	XG5838 	(WX53,WX1004,CRC_OUT_9_30);
	and 	XG5839 	(WX67,WX1004,CRC_OUT_9_29);
	and 	XG5840 	(WX81,WX1004,CRC_OUT_9_28);
	and 	XG5841 	(WX95,WX1004,CRC_OUT_9_27);
	and 	XG5842 	(WX109,WX1004,CRC_OUT_9_26);
	and 	XG5843 	(WX123,WX1004,CRC_OUT_9_25);
	and 	XG5844 	(WX137,WX1004,CRC_OUT_9_24);
	and 	XG5845 	(WX151,WX1004,CRC_OUT_9_23);
	and 	XG5846 	(WX165,WX1004,CRC_OUT_9_22);
	and 	XG5847 	(WX179,WX1004,CRC_OUT_9_21);
	and 	XG5848 	(WX193,WX1004,CRC_OUT_9_20);
	and 	XG5849 	(WX207,WX1004,CRC_OUT_9_19);
	and 	XG5850 	(WX221,WX1004,CRC_OUT_9_18);
	and 	XG5851 	(WX235,WX1004,CRC_OUT_9_17);
	and 	XG5852 	(WX249,WX1004,CRC_OUT_9_16);
	and 	XG5853 	(WX263,WX1004,CRC_OUT_9_15);
	and 	XG5854 	(WX277,WX1004,CRC_OUT_9_14);
	and 	XG5855 	(WX291,WX1004,CRC_OUT_9_13);
	and 	XG5856 	(WX305,WX1004,CRC_OUT_9_12);
	and 	XG5857 	(WX319,WX1004,CRC_OUT_9_11);
	and 	XG5858 	(WX333,WX1004,CRC_OUT_9_10);
	and 	XG5859 	(WX347,WX1004,CRC_OUT_9_9);
	and 	XG5860 	(WX361,WX1004,CRC_OUT_9_8);
	and 	XG5861 	(WX375,WX1004,CRC_OUT_9_7);
	and 	XG5862 	(WX389,WX1004,CRC_OUT_9_6);
	and 	XG5863 	(WX403,WX1004,CRC_OUT_9_5);
	and 	XG5864 	(WX417,WX1004,CRC_OUT_9_4);
	and 	XG5865 	(WX431,WX1004,CRC_OUT_9_3);
	and 	XG5866 	(WX445,WX1004,CRC_OUT_9_2);
	and 	XG5867 	(WX459,WX1004,CRC_OUT_9_1);
	and 	XG5868 	(WX473,WX1004,CRC_OUT_9_0);
	and 	XG5869 	(WX10890,RESET,WX10827);
	and 	XG5870 	(WX9597,RESET,WX9534);
	and 	XG5871 	(WX8304,RESET,WX8241);
	and 	XG5872 	(WX7011,RESET,WX6948);
	and 	XG5873 	(WX5718,RESET,WX5655);
	and 	XG5874 	(WX4425,RESET,WX4362);
	and 	XG5875 	(WX3132,RESET,WX3069);
	and 	XG5876 	(WX1839,RESET,WX1776);
	and 	XG5877 	(WX546,RESET,WX483);
	nand 	XG5878 	(II3710,CRC_OUT_9_0,WX642);
	nand 	XG5879 	(II3703,CRC_OUT_9_1,WX641);
	nand 	XG5880 	(II3696,CRC_OUT_9_2,WX640);
	nand 	XG5881 	(II3689,CRC_OUT_9_4,WX638);
	nand 	XG5882 	(II3682,CRC_OUT_9_5,WX637);
	nand 	XG5883 	(II3675,CRC_OUT_9_6,WX636);
	nand 	XG5884 	(II3668,CRC_OUT_9_7,WX635);
	nand 	XG5885 	(II3661,CRC_OUT_9_8,WX634);
	nand 	XG5886 	(II3654,CRC_OUT_9_9,WX633);
	nand 	XG5887 	(II3647,CRC_OUT_9_11,WX631);
	nand 	XG5888 	(II3640,CRC_OUT_9_12,WX630);
	nand 	XG5889 	(II3633,CRC_OUT_9_13,WX629);
	nand 	XG5890 	(II3626,CRC_OUT_9_14,WX628);
	nand 	XG5891 	(II3619,CRC_OUT_9_16,WX626);
	nand 	XG5892 	(II3612,CRC_OUT_9_17,WX625);
	nand 	XG5893 	(II3605,CRC_OUT_9_18,WX624);
	nand 	XG5894 	(II3598,CRC_OUT_9_19,WX623);
	nand 	XG5895 	(II3591,CRC_OUT_9_20,WX622);
	nand 	XG5896 	(II3584,CRC_OUT_9_21,WX621);
	nand 	XG5897 	(II3577,CRC_OUT_9_22,WX620);
	nand 	XG5898 	(II3570,CRC_OUT_9_23,WX619);
	nand 	XG5899 	(II3563,CRC_OUT_9_24,WX618);
	nand 	XG5900 	(II3556,CRC_OUT_9_25,WX617);
	nand 	XG5901 	(II3549,CRC_OUT_9_26,WX616);
	nand 	XG5902 	(II3542,CRC_OUT_9_27,WX615);
	nand 	XG5903 	(II3535,CRC_OUT_9_28,WX614);
	nand 	XG5904 	(II3528,CRC_OUT_9_29,WX613);
	nand 	XG5905 	(II3521,CRC_OUT_9_30,WX612);
	nand 	XG5906 	(II3514,CRC_OUT_9_31,WX643);
	nand 	XG5907 	(II3500,CRC_OUT_9_31,WX639);
	nand 	XG5908 	(II3485,CRC_OUT_9_31,WX632);
	nand 	XG5909 	(II3470,CRC_OUT_9_31,WX627);
	nand 	XG5910 	(II7715,CRC_OUT_8_0,WX1935);
	nand 	XG5911 	(II7708,CRC_OUT_8_1,WX1934);
	nand 	XG5912 	(II7701,CRC_OUT_8_2,WX1933);
	nand 	XG5913 	(II7694,CRC_OUT_8_4,WX1931);
	nand 	XG5914 	(II7687,CRC_OUT_8_5,WX1930);
	nand 	XG5915 	(II7680,CRC_OUT_8_6,WX1929);
	nand 	XG5916 	(II7673,CRC_OUT_8_7,WX1928);
	nand 	XG5917 	(II7666,CRC_OUT_8_8,WX1927);
	nand 	XG5918 	(II7659,CRC_OUT_8_9,WX1926);
	nand 	XG5919 	(II7652,CRC_OUT_8_11,WX1924);
	nand 	XG5920 	(II7645,CRC_OUT_8_12,WX1923);
	nand 	XG5921 	(II7638,CRC_OUT_8_13,WX1922);
	nand 	XG5922 	(II7631,CRC_OUT_8_14,WX1921);
	nand 	XG5923 	(II7624,CRC_OUT_8_16,WX1919);
	nand 	XG5924 	(II7617,CRC_OUT_8_17,WX1918);
	nand 	XG5925 	(II7610,CRC_OUT_8_18,WX1917);
	nand 	XG5926 	(II7603,CRC_OUT_8_19,WX1916);
	nand 	XG5927 	(II7596,CRC_OUT_8_20,WX1915);
	nand 	XG5928 	(II7589,CRC_OUT_8_21,WX1914);
	nand 	XG5929 	(II7582,CRC_OUT_8_22,WX1913);
	nand 	XG5930 	(II7575,CRC_OUT_8_23,WX1912);
	nand 	XG5931 	(II7568,CRC_OUT_8_24,WX1911);
	nand 	XG5932 	(II7561,CRC_OUT_8_25,WX1910);
	nand 	XG5933 	(II7554,CRC_OUT_8_26,WX1909);
	nand 	XG5934 	(II7547,CRC_OUT_8_27,WX1908);
	nand 	XG5935 	(II7540,CRC_OUT_8_28,WX1907);
	nand 	XG5936 	(II7533,CRC_OUT_8_29,WX1906);
	nand 	XG5937 	(II7526,CRC_OUT_8_30,WX1905);
	nand 	XG5938 	(II7519,CRC_OUT_8_31,WX1936);
	nand 	XG5939 	(II7505,CRC_OUT_8_31,WX1932);
	nand 	XG5940 	(II7490,CRC_OUT_8_31,WX1925);
	nand 	XG5941 	(II7475,CRC_OUT_8_31,WX1920);
	nand 	XG5942 	(II11720,CRC_OUT_7_0,WX3228);
	nand 	XG5943 	(II11713,CRC_OUT_7_1,WX3227);
	nand 	XG5944 	(II11706,CRC_OUT_7_2,WX3226);
	nand 	XG5945 	(II11699,CRC_OUT_7_4,WX3224);
	nand 	XG5946 	(II11692,CRC_OUT_7_5,WX3223);
	nand 	XG5947 	(II11685,CRC_OUT_7_6,WX3222);
	nand 	XG5948 	(II11678,CRC_OUT_7_7,WX3221);
	nand 	XG5949 	(II11671,CRC_OUT_7_8,WX3220);
	nand 	XG5950 	(II11664,CRC_OUT_7_9,WX3219);
	nand 	XG5951 	(II11657,CRC_OUT_7_11,WX3217);
	nand 	XG5952 	(II11650,CRC_OUT_7_12,WX3216);
	nand 	XG5953 	(II11643,CRC_OUT_7_13,WX3215);
	nand 	XG5954 	(II11636,CRC_OUT_7_14,WX3214);
	nand 	XG5955 	(II11629,CRC_OUT_7_16,WX3212);
	nand 	XG5956 	(II11622,CRC_OUT_7_17,WX3211);
	nand 	XG5957 	(II11615,CRC_OUT_7_18,WX3210);
	nand 	XG5958 	(II11608,CRC_OUT_7_19,WX3209);
	nand 	XG5959 	(II11601,CRC_OUT_7_20,WX3208);
	nand 	XG5960 	(II11594,CRC_OUT_7_21,WX3207);
	nand 	XG5961 	(II11587,CRC_OUT_7_22,WX3206);
	nand 	XG5962 	(II11580,CRC_OUT_7_23,WX3205);
	nand 	XG5963 	(II11573,CRC_OUT_7_24,WX3204);
	nand 	XG5964 	(II11566,CRC_OUT_7_25,WX3203);
	nand 	XG5965 	(II11559,CRC_OUT_7_26,WX3202);
	nand 	XG5966 	(II11552,CRC_OUT_7_27,WX3201);
	nand 	XG5967 	(II11545,CRC_OUT_7_28,WX3200);
	nand 	XG5968 	(II11538,CRC_OUT_7_29,WX3199);
	nand 	XG5969 	(II11531,CRC_OUT_7_30,WX3198);
	nand 	XG5970 	(II11524,CRC_OUT_7_31,WX3229);
	nand 	XG5971 	(II11510,CRC_OUT_7_31,WX3225);
	nand 	XG5972 	(II11495,CRC_OUT_7_31,WX3218);
	nand 	XG5973 	(II11480,CRC_OUT_7_31,WX3213);
	nand 	XG5974 	(II15725,CRC_OUT_6_0,WX4521);
	nand 	XG5975 	(II15718,CRC_OUT_6_1,WX4520);
	nand 	XG5976 	(II15711,CRC_OUT_6_2,WX4519);
	nand 	XG5977 	(II15704,CRC_OUT_6_4,WX4517);
	nand 	XG5978 	(II15697,CRC_OUT_6_5,WX4516);
	nand 	XG5979 	(II15690,CRC_OUT_6_6,WX4515);
	nand 	XG5980 	(II15683,CRC_OUT_6_7,WX4514);
	nand 	XG5981 	(II15676,CRC_OUT_6_8,WX4513);
	nand 	XG5982 	(II15669,CRC_OUT_6_9,WX4512);
	nand 	XG5983 	(II15662,CRC_OUT_6_11,WX4510);
	nand 	XG5984 	(II15655,CRC_OUT_6_12,WX4509);
	nand 	XG5985 	(II15648,CRC_OUT_6_13,WX4508);
	nand 	XG5986 	(II15641,CRC_OUT_6_14,WX4507);
	nand 	XG5987 	(II15634,CRC_OUT_6_16,WX4505);
	nand 	XG5988 	(II15627,CRC_OUT_6_17,WX4504);
	nand 	XG5989 	(II15620,CRC_OUT_6_18,WX4503);
	nand 	XG5990 	(II15613,CRC_OUT_6_19,WX4502);
	nand 	XG5991 	(II15606,CRC_OUT_6_20,WX4501);
	nand 	XG5992 	(II15599,CRC_OUT_6_21,WX4500);
	nand 	XG5993 	(II15592,CRC_OUT_6_22,WX4499);
	nand 	XG5994 	(II15585,CRC_OUT_6_23,WX4498);
	nand 	XG5995 	(II15578,CRC_OUT_6_24,WX4497);
	nand 	XG5996 	(II15571,CRC_OUT_6_25,WX4496);
	nand 	XG5997 	(II15564,CRC_OUT_6_26,WX4495);
	nand 	XG5998 	(II15557,CRC_OUT_6_27,WX4494);
	nand 	XG5999 	(II15550,CRC_OUT_6_28,WX4493);
	nand 	XG6000 	(II15543,CRC_OUT_6_29,WX4492);
	nand 	XG6001 	(II15536,CRC_OUT_6_30,WX4491);
	nand 	XG6002 	(II15529,CRC_OUT_6_31,WX4522);
	nand 	XG6003 	(II15515,CRC_OUT_6_31,WX4518);
	nand 	XG6004 	(II15500,CRC_OUT_6_31,WX4511);
	nand 	XG6005 	(II15485,CRC_OUT_6_31,WX4506);
	nand 	XG6006 	(II19730,CRC_OUT_5_0,WX5814);
	nand 	XG6007 	(II19723,CRC_OUT_5_1,WX5813);
	nand 	XG6008 	(II19716,CRC_OUT_5_2,WX5812);
	nand 	XG6009 	(II19709,CRC_OUT_5_4,WX5810);
	nand 	XG6010 	(II19702,CRC_OUT_5_5,WX5809);
	nand 	XG6011 	(II19695,CRC_OUT_5_6,WX5808);
	nand 	XG6012 	(II19688,CRC_OUT_5_7,WX5807);
	nand 	XG6013 	(II19681,CRC_OUT_5_8,WX5806);
	nand 	XG6014 	(II19674,CRC_OUT_5_9,WX5805);
	nand 	XG6015 	(II19667,CRC_OUT_5_11,WX5803);
	nand 	XG6016 	(II19660,CRC_OUT_5_12,WX5802);
	nand 	XG6017 	(II19653,CRC_OUT_5_13,WX5801);
	nand 	XG6018 	(II19646,CRC_OUT_5_14,WX5800);
	nand 	XG6019 	(II19639,CRC_OUT_5_16,WX5798);
	nand 	XG6020 	(II19632,CRC_OUT_5_17,WX5797);
	nand 	XG6021 	(II19625,CRC_OUT_5_18,WX5796);
	nand 	XG6022 	(II19618,CRC_OUT_5_19,WX5795);
	nand 	XG6023 	(II19611,CRC_OUT_5_20,WX5794);
	nand 	XG6024 	(II19604,CRC_OUT_5_21,WX5793);
	nand 	XG6025 	(II19597,CRC_OUT_5_22,WX5792);
	nand 	XG6026 	(II19590,CRC_OUT_5_23,WX5791);
	nand 	XG6027 	(II19583,CRC_OUT_5_24,WX5790);
	nand 	XG6028 	(II19576,CRC_OUT_5_25,WX5789);
	nand 	XG6029 	(II19569,CRC_OUT_5_26,WX5788);
	nand 	XG6030 	(II19562,CRC_OUT_5_27,WX5787);
	nand 	XG6031 	(II19555,CRC_OUT_5_28,WX5786);
	nand 	XG6032 	(II19548,CRC_OUT_5_29,WX5785);
	nand 	XG6033 	(II19541,CRC_OUT_5_30,WX5784);
	nand 	XG6034 	(II19534,CRC_OUT_5_31,WX5815);
	nand 	XG6035 	(II19520,CRC_OUT_5_31,WX5811);
	nand 	XG6036 	(II19505,CRC_OUT_5_31,WX5804);
	nand 	XG6037 	(II19490,CRC_OUT_5_31,WX5799);
	nand 	XG6038 	(II23735,CRC_OUT_4_0,WX7107);
	nand 	XG6039 	(II23728,CRC_OUT_4_1,WX7106);
	nand 	XG6040 	(II23721,CRC_OUT_4_2,WX7105);
	nand 	XG6041 	(II23714,CRC_OUT_4_4,WX7103);
	nand 	XG6042 	(II23707,CRC_OUT_4_5,WX7102);
	nand 	XG6043 	(II23700,CRC_OUT_4_6,WX7101);
	nand 	XG6044 	(II23693,CRC_OUT_4_7,WX7100);
	nand 	XG6045 	(II23686,CRC_OUT_4_8,WX7099);
	nand 	XG6046 	(II23679,CRC_OUT_4_9,WX7098);
	nand 	XG6047 	(II23672,CRC_OUT_4_11,WX7096);
	nand 	XG6048 	(II23665,CRC_OUT_4_12,WX7095);
	nand 	XG6049 	(II23658,CRC_OUT_4_13,WX7094);
	nand 	XG6050 	(II23651,CRC_OUT_4_14,WX7093);
	nand 	XG6051 	(II23644,CRC_OUT_4_16,WX7091);
	nand 	XG6052 	(II23637,CRC_OUT_4_17,WX7090);
	nand 	XG6053 	(II23630,CRC_OUT_4_18,WX7089);
	nand 	XG6054 	(II23623,CRC_OUT_4_19,WX7088);
	nand 	XG6055 	(II23616,CRC_OUT_4_20,WX7087);
	nand 	XG6056 	(II23609,CRC_OUT_4_21,WX7086);
	nand 	XG6057 	(II23602,CRC_OUT_4_22,WX7085);
	nand 	XG6058 	(II23595,CRC_OUT_4_23,WX7084);
	nand 	XG6059 	(II23588,CRC_OUT_4_24,WX7083);
	nand 	XG6060 	(II23581,CRC_OUT_4_25,WX7082);
	nand 	XG6061 	(II23574,CRC_OUT_4_26,WX7081);
	nand 	XG6062 	(II23567,CRC_OUT_4_27,WX7080);
	nand 	XG6063 	(II23560,CRC_OUT_4_28,WX7079);
	nand 	XG6064 	(II23553,CRC_OUT_4_29,WX7078);
	nand 	XG6065 	(II23546,CRC_OUT_4_30,WX7077);
	nand 	XG6066 	(II23539,CRC_OUT_4_31,WX7108);
	nand 	XG6067 	(II23525,CRC_OUT_4_31,WX7104);
	nand 	XG6068 	(II23510,CRC_OUT_4_31,WX7097);
	nand 	XG6069 	(II23495,CRC_OUT_4_31,WX7092);
	nand 	XG6070 	(II27740,CRC_OUT_3_0,WX8400);
	nand 	XG6071 	(II27733,CRC_OUT_3_1,WX8399);
	nand 	XG6072 	(II27726,CRC_OUT_3_2,WX8398);
	nand 	XG6073 	(II27719,CRC_OUT_3_4,WX8396);
	nand 	XG6074 	(II27712,CRC_OUT_3_5,WX8395);
	nand 	XG6075 	(II27705,CRC_OUT_3_6,WX8394);
	nand 	XG6076 	(II27698,CRC_OUT_3_7,WX8393);
	nand 	XG6077 	(II27691,CRC_OUT_3_8,WX8392);
	nand 	XG6078 	(II27684,CRC_OUT_3_9,WX8391);
	nand 	XG6079 	(II27677,CRC_OUT_3_11,WX8389);
	nand 	XG6080 	(II27670,CRC_OUT_3_12,WX8388);
	nand 	XG6081 	(II27663,CRC_OUT_3_13,WX8387);
	nand 	XG6082 	(II27656,CRC_OUT_3_14,WX8386);
	nand 	XG6083 	(II27649,CRC_OUT_3_16,WX8384);
	nand 	XG6084 	(II27642,CRC_OUT_3_17,WX8383);
	nand 	XG6085 	(II27635,CRC_OUT_3_18,WX8382);
	nand 	XG6086 	(II27628,CRC_OUT_3_19,WX8381);
	nand 	XG6087 	(II27621,CRC_OUT_3_20,WX8380);
	nand 	XG6088 	(II27614,CRC_OUT_3_21,WX8379);
	nand 	XG6089 	(II27607,CRC_OUT_3_22,WX8378);
	nand 	XG6090 	(II27600,CRC_OUT_3_23,WX8377);
	nand 	XG6091 	(II27593,CRC_OUT_3_24,WX8376);
	nand 	XG6092 	(II27586,CRC_OUT_3_25,WX8375);
	nand 	XG6093 	(II27579,CRC_OUT_3_26,WX8374);
	nand 	XG6094 	(II27572,CRC_OUT_3_27,WX8373);
	nand 	XG6095 	(II27565,CRC_OUT_3_28,WX8372);
	nand 	XG6096 	(II27558,CRC_OUT_3_29,WX8371);
	nand 	XG6097 	(II27551,CRC_OUT_3_30,WX8370);
	nand 	XG6098 	(II27544,CRC_OUT_3_31,WX8401);
	nand 	XG6099 	(II27530,CRC_OUT_3_31,WX8397);
	nand 	XG6100 	(II27515,CRC_OUT_3_31,WX8390);
	nand 	XG6101 	(II27500,CRC_OUT_3_31,WX8385);
	nand 	XG6102 	(II31745,CRC_OUT_2_0,WX9693);
	nand 	XG6103 	(II31738,CRC_OUT_2_1,WX9692);
	nand 	XG6104 	(II31731,CRC_OUT_2_2,WX9691);
	nand 	XG6105 	(II31724,CRC_OUT_2_4,WX9689);
	nand 	XG6106 	(II31717,CRC_OUT_2_5,WX9688);
	nand 	XG6107 	(II31710,CRC_OUT_2_6,WX9687);
	nand 	XG6108 	(II31703,CRC_OUT_2_7,WX9686);
	nand 	XG6109 	(II31696,CRC_OUT_2_8,WX9685);
	nand 	XG6110 	(II31689,CRC_OUT_2_9,WX9684);
	nand 	XG6111 	(II31682,CRC_OUT_2_11,WX9682);
	nand 	XG6112 	(II31675,CRC_OUT_2_12,WX9681);
	nand 	XG6113 	(II31668,CRC_OUT_2_13,WX9680);
	nand 	XG6114 	(II31661,CRC_OUT_2_14,WX9679);
	nand 	XG6115 	(II31654,CRC_OUT_2_16,WX9677);
	nand 	XG6116 	(II31647,CRC_OUT_2_17,WX9676);
	nand 	XG6117 	(II31640,CRC_OUT_2_18,WX9675);
	nand 	XG6118 	(II31633,CRC_OUT_2_19,WX9674);
	nand 	XG6119 	(II31626,CRC_OUT_2_20,WX9673);
	nand 	XG6120 	(II31619,CRC_OUT_2_21,WX9672);
	nand 	XG6121 	(II31612,CRC_OUT_2_22,WX9671);
	nand 	XG6122 	(II31605,CRC_OUT_2_23,WX9670);
	nand 	XG6123 	(II31598,CRC_OUT_2_24,WX9669);
	nand 	XG6124 	(II31591,CRC_OUT_2_25,WX9668);
	nand 	XG6125 	(II31584,CRC_OUT_2_26,WX9667);
	nand 	XG6126 	(II31577,CRC_OUT_2_27,WX9666);
	nand 	XG6127 	(II31570,CRC_OUT_2_28,WX9665);
	nand 	XG6128 	(II31563,CRC_OUT_2_29,WX9664);
	nand 	XG6129 	(II31556,CRC_OUT_2_30,WX9663);
	nand 	XG6130 	(II31549,CRC_OUT_2_31,WX9694);
	nand 	XG6131 	(II31535,CRC_OUT_2_31,WX9690);
	nand 	XG6132 	(II31520,CRC_OUT_2_31,WX9683);
	nand 	XG6133 	(II31505,CRC_OUT_2_31,WX9678);
	nand 	XG6134 	(II35750,CRC_OUT_1_0,WX10986);
	nand 	XG6135 	(II35743,CRC_OUT_1_1,WX10985);
	nand 	XG6136 	(II35736,CRC_OUT_1_2,WX10984);
	nand 	XG6137 	(II35729,CRC_OUT_1_4,WX10982);
	nand 	XG6138 	(II35722,CRC_OUT_1_5,WX10981);
	nand 	XG6139 	(II35715,CRC_OUT_1_6,WX10980);
	nand 	XG6140 	(II35708,CRC_OUT_1_7,WX10979);
	nand 	XG6141 	(II35701,CRC_OUT_1_8,WX10978);
	nand 	XG6142 	(II35694,CRC_OUT_1_9,WX10977);
	nand 	XG6143 	(II35687,CRC_OUT_1_11,WX10975);
	nand 	XG6144 	(II35680,CRC_OUT_1_12,WX10974);
	nand 	XG6145 	(II35673,CRC_OUT_1_13,WX10973);
	nand 	XG6146 	(II35666,CRC_OUT_1_14,WX10972);
	nand 	XG6147 	(II35659,CRC_OUT_1_16,WX10970);
	nand 	XG6148 	(II35652,CRC_OUT_1_17,WX10969);
	nand 	XG6149 	(II35645,CRC_OUT_1_18,WX10968);
	nand 	XG6150 	(II35638,CRC_OUT_1_19,WX10967);
	nand 	XG6151 	(II35631,CRC_OUT_1_20,WX10966);
	nand 	XG6152 	(II35624,CRC_OUT_1_21,WX10965);
	nand 	XG6153 	(II35617,CRC_OUT_1_22,WX10964);
	nand 	XG6154 	(II35610,CRC_OUT_1_23,WX10963);
	nand 	XG6155 	(II35603,CRC_OUT_1_24,WX10962);
	nand 	XG6156 	(II35596,CRC_OUT_1_25,WX10961);
	nand 	XG6157 	(II35589,CRC_OUT_1_26,WX10960);
	nand 	XG6158 	(II35582,CRC_OUT_1_27,WX10959);
	nand 	XG6159 	(II35575,CRC_OUT_1_28,WX10958);
	nand 	XG6160 	(II35568,CRC_OUT_1_29,WX10957);
	nand 	XG6161 	(II35561,CRC_OUT_1_30,WX10956);
	nand 	XG6162 	(II35554,CRC_OUT_1_31,WX10987);
	nand 	XG6163 	(II35540,CRC_OUT_1_31,WX10983);
	nand 	XG6164 	(II35525,CRC_OUT_1_31,WX10976);
	nand 	XG6165 	(II35510,CRC_OUT_1_31,WX10971);
	nand 	XG6166 	(II2004,II2003,WX773);
	nand 	XG6167 	(II2035,II2034,WX775);
	nand 	XG6168 	(II2066,II2065,WX777);
	nand 	XG6169 	(II2097,II2096,WX779);
	nand 	XG6170 	(II2128,II2127,WX781);
	nand 	XG6171 	(II2159,II2158,WX783);
	nand 	XG6172 	(II2190,II2189,WX785);
	nand 	XG6173 	(II2221,II2220,WX787);
	nand 	XG6174 	(II2252,II2251,WX789);
	nand 	XG6175 	(II2283,II2282,WX791);
	nand 	XG6176 	(II2314,II2313,WX793);
	nand 	XG6177 	(II2345,II2344,WX795);
	nand 	XG6178 	(II2376,II2375,WX797);
	nand 	XG6179 	(II2407,II2406,WX799);
	nand 	XG6180 	(II2438,II2437,WX801);
	nand 	XG6181 	(II2469,II2468,WX803);
	nand 	XG6182 	(II2500,II2499,WX805);
	nand 	XG6183 	(II2531,II2530,WX807);
	nand 	XG6184 	(II2562,II2561,WX809);
	nand 	XG6185 	(II2593,II2592,WX811);
	nand 	XG6186 	(II2624,II2623,WX813);
	nand 	XG6187 	(II2655,II2654,WX815);
	nand 	XG6188 	(II2686,II2685,WX817);
	nand 	XG6189 	(II2717,II2716,WX819);
	nand 	XG6190 	(II2748,II2747,WX821);
	nand 	XG6191 	(II2779,II2778,WX823);
	nand 	XG6192 	(II2810,II2809,WX825);
	nand 	XG6193 	(II2841,II2840,WX827);
	nand 	XG6194 	(II2872,II2871,WX829);
	nand 	XG6195 	(II2903,II2902,WX831);
	nand 	XG6196 	(II2934,II2933,WX833);
	nand 	XG6197 	(II2965,II2964,WX835);
	nand 	XG6198 	(II6009,II6008,WX2066);
	nand 	XG6199 	(II6040,II6039,WX2068);
	nand 	XG6200 	(II6071,II6070,WX2070);
	nand 	XG6201 	(II6102,II6101,WX2072);
	nand 	XG6202 	(II6133,II6132,WX2074);
	nand 	XG6203 	(II6164,II6163,WX2076);
	nand 	XG6204 	(II6195,II6194,WX2078);
	nand 	XG6205 	(II6226,II6225,WX2080);
	nand 	XG6206 	(II6257,II6256,WX2082);
	nand 	XG6207 	(II6288,II6287,WX2084);
	nand 	XG6208 	(II6319,II6318,WX2086);
	nand 	XG6209 	(II6350,II6349,WX2088);
	nand 	XG6210 	(II6381,II6380,WX2090);
	nand 	XG6211 	(II6412,II6411,WX2092);
	nand 	XG6212 	(II6443,II6442,WX2094);
	nand 	XG6213 	(II6474,II6473,WX2096);
	nand 	XG6214 	(II6505,II6504,WX2098);
	nand 	XG6215 	(II6536,II6535,WX2100);
	nand 	XG6216 	(II6567,II6566,WX2102);
	nand 	XG6217 	(II6598,II6597,WX2104);
	nand 	XG6218 	(II6629,II6628,WX2106);
	nand 	XG6219 	(II6660,II6659,WX2108);
	nand 	XG6220 	(II6691,II6690,WX2110);
	nand 	XG6221 	(II6722,II6721,WX2112);
	nand 	XG6222 	(II6753,II6752,WX2114);
	nand 	XG6223 	(II6784,II6783,WX2116);
	nand 	XG6224 	(II6815,II6814,WX2118);
	nand 	XG6225 	(II6846,II6845,WX2120);
	nand 	XG6226 	(II6877,II6876,WX2122);
	nand 	XG6227 	(II6908,II6907,WX2124);
	nand 	XG6228 	(II6939,II6938,WX2126);
	nand 	XG6229 	(II6970,II6969,WX2128);
	nand 	XG6230 	(II10014,II10013,WX3359);
	nand 	XG6231 	(II10045,II10044,WX3361);
	nand 	XG6232 	(II10076,II10075,WX3363);
	nand 	XG6233 	(II10107,II10106,WX3365);
	nand 	XG6234 	(II10138,II10137,WX3367);
	nand 	XG6235 	(II10169,II10168,WX3369);
	nand 	XG6236 	(II10200,II10199,WX3371);
	nand 	XG6237 	(II10231,II10230,WX3373);
	nand 	XG6238 	(II10262,II10261,WX3375);
	nand 	XG6239 	(II10293,II10292,WX3377);
	nand 	XG6240 	(II10324,II10323,WX3379);
	nand 	XG6241 	(II10355,II10354,WX3381);
	nand 	XG6242 	(II10386,II10385,WX3383);
	nand 	XG6243 	(II10417,II10416,WX3385);
	nand 	XG6244 	(II10448,II10447,WX3387);
	nand 	XG6245 	(II10479,II10478,WX3389);
	nand 	XG6246 	(II10510,II10509,WX3391);
	nand 	XG6247 	(II10541,II10540,WX3393);
	nand 	XG6248 	(II10572,II10571,WX3395);
	nand 	XG6249 	(II10603,II10602,WX3397);
	nand 	XG6250 	(II10634,II10633,WX3399);
	nand 	XG6251 	(II10665,II10664,WX3401);
	nand 	XG6252 	(II10696,II10695,WX3403);
	nand 	XG6253 	(II10727,II10726,WX3405);
	nand 	XG6254 	(II10758,II10757,WX3407);
	nand 	XG6255 	(II10789,II10788,WX3409);
	nand 	XG6256 	(II10820,II10819,WX3411);
	nand 	XG6257 	(II10851,II10850,WX3413);
	nand 	XG6258 	(II10882,II10881,WX3415);
	nand 	XG6259 	(II10913,II10912,WX3417);
	nand 	XG6260 	(II10944,II10943,WX3419);
	nand 	XG6261 	(II10975,II10974,WX3421);
	nand 	XG6262 	(II14019,II14018,WX4652);
	nand 	XG6263 	(II14050,II14049,WX4654);
	nand 	XG6264 	(II14081,II14080,WX4656);
	nand 	XG6265 	(II14112,II14111,WX4658);
	nand 	XG6266 	(II14143,II14142,WX4660);
	nand 	XG6267 	(II14174,II14173,WX4662);
	nand 	XG6268 	(II14205,II14204,WX4664);
	nand 	XG6269 	(II14236,II14235,WX4666);
	nand 	XG6270 	(II14267,II14266,WX4668);
	nand 	XG6271 	(II14298,II14297,WX4670);
	nand 	XG6272 	(II14329,II14328,WX4672);
	nand 	XG6273 	(II14360,II14359,WX4674);
	nand 	XG6274 	(II14391,II14390,WX4676);
	nand 	XG6275 	(II14422,II14421,WX4678);
	nand 	XG6276 	(II14453,II14452,WX4680);
	nand 	XG6277 	(II14484,II14483,WX4682);
	nand 	XG6278 	(II14515,II14514,WX4684);
	nand 	XG6279 	(II14546,II14545,WX4686);
	nand 	XG6280 	(II14577,II14576,WX4688);
	nand 	XG6281 	(II14608,II14607,WX4690);
	nand 	XG6282 	(II14639,II14638,WX4692);
	nand 	XG6283 	(II14670,II14669,WX4694);
	nand 	XG6284 	(II14701,II14700,WX4696);
	nand 	XG6285 	(II14732,II14731,WX4698);
	nand 	XG6286 	(II14763,II14762,WX4700);
	nand 	XG6287 	(II14794,II14793,WX4702);
	nand 	XG6288 	(II14825,II14824,WX4704);
	nand 	XG6289 	(II14856,II14855,WX4706);
	nand 	XG6290 	(II14887,II14886,WX4708);
	nand 	XG6291 	(II14918,II14917,WX4710);
	nand 	XG6292 	(II14949,II14948,WX4712);
	nand 	XG6293 	(II14980,II14979,WX4714);
	nand 	XG6294 	(II18024,II18023,WX5945);
	nand 	XG6295 	(II18055,II18054,WX5947);
	nand 	XG6296 	(II18086,II18085,WX5949);
	nand 	XG6297 	(II18117,II18116,WX5951);
	nand 	XG6298 	(II18148,II18147,WX5953);
	nand 	XG6299 	(II18179,II18178,WX5955);
	nand 	XG6300 	(II18210,II18209,WX5957);
	nand 	XG6301 	(II18241,II18240,WX5959);
	nand 	XG6302 	(II18272,II18271,WX5961);
	nand 	XG6303 	(II18303,II18302,WX5963);
	nand 	XG6304 	(II18334,II18333,WX5965);
	nand 	XG6305 	(II18365,II18364,WX5967);
	nand 	XG6306 	(II18396,II18395,WX5969);
	nand 	XG6307 	(II18427,II18426,WX5971);
	nand 	XG6308 	(II18458,II18457,WX5973);
	nand 	XG6309 	(II18489,II18488,WX5975);
	nand 	XG6310 	(II18520,II18519,WX5977);
	nand 	XG6311 	(II18551,II18550,WX5979);
	nand 	XG6312 	(II18582,II18581,WX5981);
	nand 	XG6313 	(II18613,II18612,WX5983);
	nand 	XG6314 	(II18644,II18643,WX5985);
	nand 	XG6315 	(II18675,II18674,WX5987);
	nand 	XG6316 	(II18706,II18705,WX5989);
	nand 	XG6317 	(II18737,II18736,WX5991);
	nand 	XG6318 	(II18768,II18767,WX5993);
	nand 	XG6319 	(II18799,II18798,WX5995);
	nand 	XG6320 	(II18830,II18829,WX5997);
	nand 	XG6321 	(II18861,II18860,WX5999);
	nand 	XG6322 	(II18892,II18891,WX6001);
	nand 	XG6323 	(II18923,II18922,WX6003);
	nand 	XG6324 	(II18954,II18953,WX6005);
	nand 	XG6325 	(II18985,II18984,WX6007);
	nand 	XG6326 	(II22029,II22028,WX7238);
	nand 	XG6327 	(II22060,II22059,WX7240);
	nand 	XG6328 	(II22091,II22090,WX7242);
	nand 	XG6329 	(II22122,II22121,WX7244);
	nand 	XG6330 	(II22153,II22152,WX7246);
	nand 	XG6331 	(II22184,II22183,WX7248);
	nand 	XG6332 	(II22215,II22214,WX7250);
	nand 	XG6333 	(II22246,II22245,WX7252);
	nand 	XG6334 	(II22277,II22276,WX7254);
	nand 	XG6335 	(II22308,II22307,WX7256);
	nand 	XG6336 	(II22339,II22338,WX7258);
	nand 	XG6337 	(II22370,II22369,WX7260);
	nand 	XG6338 	(II22401,II22400,WX7262);
	nand 	XG6339 	(II22432,II22431,WX7264);
	nand 	XG6340 	(II22463,II22462,WX7266);
	nand 	XG6341 	(II22494,II22493,WX7268);
	nand 	XG6342 	(II22525,II22524,WX7270);
	nand 	XG6343 	(II22556,II22555,WX7272);
	nand 	XG6344 	(II22587,II22586,WX7274);
	nand 	XG6345 	(II22618,II22617,WX7276);
	nand 	XG6346 	(II22649,II22648,WX7278);
	nand 	XG6347 	(II22680,II22679,WX7280);
	nand 	XG6348 	(II22711,II22710,WX7282);
	nand 	XG6349 	(II22742,II22741,WX7284);
	nand 	XG6350 	(II22773,II22772,WX7286);
	nand 	XG6351 	(II22804,II22803,WX7288);
	nand 	XG6352 	(II22835,II22834,WX7290);
	nand 	XG6353 	(II22866,II22865,WX7292);
	nand 	XG6354 	(II22897,II22896,WX7294);
	nand 	XG6355 	(II22928,II22927,WX7296);
	nand 	XG6356 	(II22959,II22958,WX7298);
	nand 	XG6357 	(II22990,II22989,WX7300);
	nand 	XG6358 	(II26034,II26033,WX8531);
	nand 	XG6359 	(II26065,II26064,WX8533);
	nand 	XG6360 	(II26096,II26095,WX8535);
	nand 	XG6361 	(II26127,II26126,WX8537);
	nand 	XG6362 	(II26158,II26157,WX8539);
	nand 	XG6363 	(II26189,II26188,WX8541);
	nand 	XG6364 	(II26220,II26219,WX8543);
	nand 	XG6365 	(II26251,II26250,WX8545);
	nand 	XG6366 	(II26282,II26281,WX8547);
	nand 	XG6367 	(II26313,II26312,WX8549);
	nand 	XG6368 	(II26344,II26343,WX8551);
	nand 	XG6369 	(II26375,II26374,WX8553);
	nand 	XG6370 	(II26406,II26405,WX8555);
	nand 	XG6371 	(II26437,II26436,WX8557);
	nand 	XG6372 	(II26468,II26467,WX8559);
	nand 	XG6373 	(II26499,II26498,WX8561);
	nand 	XG6374 	(II26530,II26529,WX8563);
	nand 	XG6375 	(II26561,II26560,WX8565);
	nand 	XG6376 	(II26592,II26591,WX8567);
	nand 	XG6377 	(II26623,II26622,WX8569);
	nand 	XG6378 	(II26654,II26653,WX8571);
	nand 	XG6379 	(II26685,II26684,WX8573);
	nand 	XG6380 	(II26716,II26715,WX8575);
	nand 	XG6381 	(II26747,II26746,WX8577);
	nand 	XG6382 	(II26778,II26777,WX8579);
	nand 	XG6383 	(II26809,II26808,WX8581);
	nand 	XG6384 	(II26840,II26839,WX8583);
	nand 	XG6385 	(II26871,II26870,WX8585);
	nand 	XG6386 	(II26902,II26901,WX8587);
	nand 	XG6387 	(II26933,II26932,WX8589);
	nand 	XG6388 	(II26964,II26963,WX8591);
	nand 	XG6389 	(II26995,II26994,WX8593);
	nand 	XG6390 	(II30039,II30038,WX9824);
	nand 	XG6391 	(II30070,II30069,WX9826);
	nand 	XG6392 	(II30101,II30100,WX9828);
	nand 	XG6393 	(II30132,II30131,WX9830);
	nand 	XG6394 	(II30163,II30162,WX9832);
	nand 	XG6395 	(II30194,II30193,WX9834);
	nand 	XG6396 	(II30225,II30224,WX9836);
	nand 	XG6397 	(II30256,II30255,WX9838);
	nand 	XG6398 	(II30287,II30286,WX9840);
	nand 	XG6399 	(II30318,II30317,WX9842);
	nand 	XG6400 	(II30349,II30348,WX9844);
	nand 	XG6401 	(II30380,II30379,WX9846);
	nand 	XG6402 	(II30411,II30410,WX9848);
	nand 	XG6403 	(II30442,II30441,WX9850);
	nand 	XG6404 	(II30473,II30472,WX9852);
	nand 	XG6405 	(II30504,II30503,WX9854);
	nand 	XG6406 	(II30535,II30534,WX9856);
	nand 	XG6407 	(II30566,II30565,WX9858);
	nand 	XG6408 	(II30597,II30596,WX9860);
	nand 	XG6409 	(II30628,II30627,WX9862);
	nand 	XG6410 	(II30659,II30658,WX9864);
	nand 	XG6411 	(II30690,II30689,WX9866);
	nand 	XG6412 	(II30721,II30720,WX9868);
	nand 	XG6413 	(II30752,II30751,WX9870);
	nand 	XG6414 	(II30783,II30782,WX9872);
	nand 	XG6415 	(II30814,II30813,WX9874);
	nand 	XG6416 	(II30845,II30844,WX9876);
	nand 	XG6417 	(II30876,II30875,WX9878);
	nand 	XG6418 	(II30907,II30906,WX9880);
	nand 	XG6419 	(II30938,II30937,WX9882);
	nand 	XG6420 	(II30969,II30968,WX9884);
	nand 	XG6421 	(II31000,II30999,WX9886);
	nand 	XG6422 	(II34044,II34043,WX11117);
	nand 	XG6423 	(II34075,II34074,WX11119);
	nand 	XG6424 	(II34106,II34105,WX11121);
	nand 	XG6425 	(II34137,II34136,WX11123);
	nand 	XG6426 	(II34168,II34167,WX11125);
	nand 	XG6427 	(II34199,II34198,WX11127);
	nand 	XG6428 	(II34230,II34229,WX11129);
	nand 	XG6429 	(II34261,II34260,WX11131);
	nand 	XG6430 	(II34292,II34291,WX11133);
	nand 	XG6431 	(II34323,II34322,WX11135);
	nand 	XG6432 	(II34354,II34353,WX11137);
	nand 	XG6433 	(II34385,II34384,WX11139);
	nand 	XG6434 	(II34416,II34415,WX11141);
	nand 	XG6435 	(II34447,II34446,WX11143);
	nand 	XG6436 	(II34478,II34477,WX11145);
	nand 	XG6437 	(II34509,II34508,WX11147);
	nand 	XG6438 	(II34540,II34539,WX11149);
	nand 	XG6439 	(II34571,II34570,WX11151);
	nand 	XG6440 	(II34602,II34601,WX11153);
	nand 	XG6441 	(II34633,II34632,WX11155);
	nand 	XG6442 	(II34664,II34663,WX11157);
	nand 	XG6443 	(II34695,II34694,WX11159);
	nand 	XG6444 	(II34726,II34725,WX11161);
	nand 	XG6445 	(II34757,II34756,WX11163);
	nand 	XG6446 	(II34788,II34787,WX11165);
	nand 	XG6447 	(II34819,II34818,WX11167);
	nand 	XG6448 	(II34850,II34849,WX11169);
	nand 	XG6449 	(II34881,II34880,WX11171);
	nand 	XG6450 	(II34912,II34911,WX11173);
	nand 	XG6451 	(II34943,II34942,WX11175);
	nand 	XG6452 	(II34974,II34973,WX11177);
	nand 	XG6453 	(II35005,II35004,WX11179);
	and 	XG6454 	(WX10384,WX10385,DATA_0_31);
	and 	XG6455 	(WX10398,WX10399,DATA_0_30);
	and 	XG6456 	(WX10412,WX10413,DATA_0_29);
	and 	XG6457 	(WX10426,WX10427,DATA_0_28);
	and 	XG6458 	(WX10440,WX10441,DATA_0_27);
	and 	XG6459 	(WX10454,WX10455,DATA_0_26);
	and 	XG6460 	(WX10468,WX10469,DATA_0_25);
	and 	XG6461 	(WX10482,WX10483,DATA_0_24);
	and 	XG6462 	(WX10496,WX10497,DATA_0_23);
	and 	XG6463 	(WX10510,WX10511,DATA_0_22);
	and 	XG6464 	(WX10524,WX10525,DATA_0_21);
	and 	XG6465 	(WX10538,WX10539,DATA_0_20);
	and 	XG6466 	(WX10552,WX10553,DATA_0_19);
	and 	XG6467 	(WX10566,WX10567,DATA_0_18);
	and 	XG6468 	(WX10580,WX10581,DATA_0_17);
	and 	XG6469 	(WX10594,WX10595,DATA_0_16);
	and 	XG6470 	(WX10608,WX10609,DATA_0_15);
	and 	XG6471 	(WX10622,WX10623,DATA_0_14);
	and 	XG6472 	(WX10636,WX10637,DATA_0_13);
	and 	XG6473 	(WX10650,WX10651,DATA_0_12);
	and 	XG6474 	(WX10664,WX10665,DATA_0_11);
	and 	XG6475 	(WX10678,WX10679,DATA_0_10);
	and 	XG6476 	(WX10692,WX10693,DATA_0_9);
	and 	XG6477 	(WX10706,WX10707,DATA_0_8);
	and 	XG6478 	(WX10720,WX10721,DATA_0_7);
	and 	XG6479 	(WX10734,WX10735,DATA_0_6);
	and 	XG6480 	(WX10748,WX10749,DATA_0_5);
	and 	XG6481 	(WX10762,WX10763,DATA_0_4);
	and 	XG6482 	(WX10776,WX10777,DATA_0_3);
	and 	XG6483 	(WX10790,WX10791,DATA_0_2);
	and 	XG6484 	(WX10804,WX10805,DATA_0_1);
	and 	XG6485 	(WX10818,WX10819,DATA_0_0);
	nand 	XG6486 	(II34494,II34493,WX11345);
	nand 	XG6487 	(II34463,II34462,WX11345);
	nand 	XG6488 	(II34432,II34431,WX11345);
	nand 	XG6489 	(II34401,II34400,WX11345);
	nand 	XG6490 	(II34370,II34369,WX11345);
	nand 	XG6491 	(II34339,II34338,WX11345);
	nand 	XG6492 	(II34308,II34307,WX11345);
	nand 	XG6493 	(II34277,II34276,WX11345);
	nand 	XG6494 	(II34246,II34245,WX11345);
	nand 	XG6495 	(II34215,II34214,WX11345);
	nand 	XG6496 	(II34184,II34183,WX11345);
	nand 	XG6497 	(II34153,II34152,WX11345);
	nand 	XG6498 	(II34122,II34121,WX11345);
	nand 	XG6499 	(II34091,II34090,WX11345);
	nand 	XG6500 	(II34060,II34059,WX11345);
	nand 	XG6501 	(II34029,II34028,WX11345);
	nand 	XG6502 	(II30489,II30488,WX10052);
	nand 	XG6503 	(II30458,II30457,WX10052);
	nand 	XG6504 	(II30427,II30426,WX10052);
	nand 	XG6505 	(II30396,II30395,WX10052);
	nand 	XG6506 	(II30365,II30364,WX10052);
	nand 	XG6507 	(II30334,II30333,WX10052);
	nand 	XG6508 	(II30303,II30302,WX10052);
	nand 	XG6509 	(II30272,II30271,WX10052);
	nand 	XG6510 	(II30241,II30240,WX10052);
	nand 	XG6511 	(II30210,II30209,WX10052);
	nand 	XG6512 	(II30179,II30178,WX10052);
	nand 	XG6513 	(II30148,II30147,WX10052);
	nand 	XG6514 	(II30117,II30116,WX10052);
	nand 	XG6515 	(II30086,II30085,WX10052);
	nand 	XG6516 	(II30055,II30054,WX10052);
	nand 	XG6517 	(II30024,II30023,WX10052);
	nand 	XG6518 	(II26484,II26483,WX8759);
	nand 	XG6519 	(II26453,II26452,WX8759);
	nand 	XG6520 	(II26422,II26421,WX8759);
	nand 	XG6521 	(II26391,II26390,WX8759);
	nand 	XG6522 	(II26360,II26359,WX8759);
	nand 	XG6523 	(II26329,II26328,WX8759);
	nand 	XG6524 	(II26298,II26297,WX8759);
	nand 	XG6525 	(II26267,II26266,WX8759);
	nand 	XG6526 	(II26236,II26235,WX8759);
	nand 	XG6527 	(II26205,II26204,WX8759);
	nand 	XG6528 	(II26174,II26173,WX8759);
	nand 	XG6529 	(II26143,II26142,WX8759);
	nand 	XG6530 	(II26112,II26111,WX8759);
	nand 	XG6531 	(II26081,II26080,WX8759);
	nand 	XG6532 	(II26050,II26049,WX8759);
	nand 	XG6533 	(II26019,II26018,WX8759);
	nand 	XG6534 	(II22479,II22478,WX7466);
	nand 	XG6535 	(II22448,II22447,WX7466);
	nand 	XG6536 	(II22417,II22416,WX7466);
	nand 	XG6537 	(II22386,II22385,WX7466);
	nand 	XG6538 	(II22355,II22354,WX7466);
	nand 	XG6539 	(II22324,II22323,WX7466);
	nand 	XG6540 	(II22293,II22292,WX7466);
	nand 	XG6541 	(II22262,II22261,WX7466);
	nand 	XG6542 	(II22231,II22230,WX7466);
	nand 	XG6543 	(II22200,II22199,WX7466);
	nand 	XG6544 	(II22169,II22168,WX7466);
	nand 	XG6545 	(II22138,II22137,WX7466);
	nand 	XG6546 	(II22107,II22106,WX7466);
	nand 	XG6547 	(II22076,II22075,WX7466);
	nand 	XG6548 	(II22045,II22044,WX7466);
	nand 	XG6549 	(II22014,II22013,WX7466);
	nand 	XG6550 	(II18474,II18473,WX6173);
	nand 	XG6551 	(II18443,II18442,WX6173);
	nand 	XG6552 	(II18412,II18411,WX6173);
	nand 	XG6553 	(II18381,II18380,WX6173);
	nand 	XG6554 	(II18350,II18349,WX6173);
	nand 	XG6555 	(II18319,II18318,WX6173);
	nand 	XG6556 	(II18288,II18287,WX6173);
	nand 	XG6557 	(II18257,II18256,WX6173);
	nand 	XG6558 	(II18226,II18225,WX6173);
	nand 	XG6559 	(II18195,II18194,WX6173);
	nand 	XG6560 	(II18164,II18163,WX6173);
	nand 	XG6561 	(II18133,II18132,WX6173);
	nand 	XG6562 	(II18102,II18101,WX6173);
	nand 	XG6563 	(II18071,II18070,WX6173);
	nand 	XG6564 	(II18040,II18039,WX6173);
	nand 	XG6565 	(II18009,II18008,WX6173);
	nand 	XG6566 	(II14469,II14468,WX4880);
	nand 	XG6567 	(II14438,II14437,WX4880);
	nand 	XG6568 	(II14407,II14406,WX4880);
	nand 	XG6569 	(II14376,II14375,WX4880);
	nand 	XG6570 	(II14345,II14344,WX4880);
	nand 	XG6571 	(II14314,II14313,WX4880);
	nand 	XG6572 	(II14283,II14282,WX4880);
	nand 	XG6573 	(II14252,II14251,WX4880);
	nand 	XG6574 	(II14221,II14220,WX4880);
	nand 	XG6575 	(II14190,II14189,WX4880);
	nand 	XG6576 	(II14159,II14158,WX4880);
	nand 	XG6577 	(II14128,II14127,WX4880);
	nand 	XG6578 	(II14097,II14096,WX4880);
	nand 	XG6579 	(II14066,II14065,WX4880);
	nand 	XG6580 	(II14035,II14034,WX4880);
	nand 	XG6581 	(II14004,II14003,WX4880);
	nand 	XG6582 	(II10464,II10463,WX3587);
	nand 	XG6583 	(II10433,II10432,WX3587);
	nand 	XG6584 	(II10402,II10401,WX3587);
	nand 	XG6585 	(II10371,II10370,WX3587);
	nand 	XG6586 	(II10340,II10339,WX3587);
	nand 	XG6587 	(II10309,II10308,WX3587);
	nand 	XG6588 	(II10278,II10277,WX3587);
	nand 	XG6589 	(II10247,II10246,WX3587);
	nand 	XG6590 	(II10216,II10215,WX3587);
	nand 	XG6591 	(II10185,II10184,WX3587);
	nand 	XG6592 	(II10154,II10153,WX3587);
	nand 	XG6593 	(II10123,II10122,WX3587);
	nand 	XG6594 	(II10092,II10091,WX3587);
	nand 	XG6595 	(II10061,II10060,WX3587);
	nand 	XG6596 	(II10030,II10029,WX3587);
	nand 	XG6597 	(II9999,II9998,WX3587);
	nand 	XG6598 	(II6459,II6458,WX2294);
	nand 	XG6599 	(II6428,II6427,WX2294);
	nand 	XG6600 	(II6397,II6396,WX2294);
	nand 	XG6601 	(II6366,II6365,WX2294);
	nand 	XG6602 	(II6335,II6334,WX2294);
	nand 	XG6603 	(II6304,II6303,WX2294);
	nand 	XG6604 	(II6273,II6272,WX2294);
	nand 	XG6605 	(II6242,II6241,WX2294);
	nand 	XG6606 	(II6211,II6210,WX2294);
	nand 	XG6607 	(II6180,II6179,WX2294);
	nand 	XG6608 	(II6149,II6148,WX2294);
	nand 	XG6609 	(II6118,II6117,WX2294);
	nand 	XG6610 	(II6087,II6086,WX2294);
	nand 	XG6611 	(II6056,II6055,WX2294);
	nand 	XG6612 	(II6025,II6024,WX2294);
	nand 	XG6613 	(II5994,II5993,WX2294);
	nand 	XG6614 	(II2454,II2453,WX1001);
	nand 	XG6615 	(II2423,II2422,WX1001);
	nand 	XG6616 	(II2392,II2391,WX1001);
	nand 	XG6617 	(II2361,II2360,WX1001);
	nand 	XG6618 	(II2330,II2329,WX1001);
	nand 	XG6619 	(II2299,II2298,WX1001);
	nand 	XG6620 	(II2268,II2267,WX1001);
	nand 	XG6621 	(II2237,II2236,WX1001);
	nand 	XG6622 	(II2206,II2205,WX1001);
	nand 	XG6623 	(II2175,II2174,WX1001);
	nand 	XG6624 	(II2144,II2143,WX1001);
	nand 	XG6625 	(II2113,II2112,WX1001);
	nand 	XG6626 	(II2082,II2081,WX1001);
	nand 	XG6627 	(II2051,II2050,WX1001);
	nand 	XG6628 	(II2020,II2019,WX1001);
	nand 	XG6629 	(II1989,II1988,WX1001);
	nand 	XG6630 	(II34990,II34989,WX11346);
	nand 	XG6631 	(II34959,II34958,WX11346);
	nand 	XG6632 	(II34928,II34927,WX11346);
	nand 	XG6633 	(II34897,II34896,WX11346);
	nand 	XG6634 	(II34866,II34865,WX11346);
	nand 	XG6635 	(II34835,II34834,WX11346);
	nand 	XG6636 	(II34804,II34803,WX11346);
	nand 	XG6637 	(II34773,II34772,WX11346);
	nand 	XG6638 	(II34742,II34741,WX11346);
	nand 	XG6639 	(II34711,II34710,WX11346);
	nand 	XG6640 	(II34680,II34679,WX11346);
	nand 	XG6641 	(II34649,II34648,WX11346);
	nand 	XG6642 	(II34618,II34617,WX11346);
	nand 	XG6643 	(II34587,II34586,WX11346);
	nand 	XG6644 	(II34556,II34555,WX11346);
	nand 	XG6645 	(II34525,II34524,WX11346);
	nand 	XG6646 	(II30985,II30984,WX10053);
	nand 	XG6647 	(II30954,II30953,WX10053);
	nand 	XG6648 	(II30923,II30922,WX10053);
	nand 	XG6649 	(II30892,II30891,WX10053);
	nand 	XG6650 	(II30861,II30860,WX10053);
	nand 	XG6651 	(II30830,II30829,WX10053);
	nand 	XG6652 	(II30799,II30798,WX10053);
	nand 	XG6653 	(II30768,II30767,WX10053);
	nand 	XG6654 	(II30737,II30736,WX10053);
	nand 	XG6655 	(II30706,II30705,WX10053);
	nand 	XG6656 	(II30675,II30674,WX10053);
	nand 	XG6657 	(II30644,II30643,WX10053);
	nand 	XG6658 	(II30613,II30612,WX10053);
	nand 	XG6659 	(II30582,II30581,WX10053);
	nand 	XG6660 	(II30551,II30550,WX10053);
	nand 	XG6661 	(II30520,II30519,WX10053);
	nand 	XG6662 	(II26980,II26979,WX8760);
	nand 	XG6663 	(II26949,II26948,WX8760);
	nand 	XG6664 	(II26918,II26917,WX8760);
	nand 	XG6665 	(II26887,II26886,WX8760);
	nand 	XG6666 	(II26856,II26855,WX8760);
	nand 	XG6667 	(II26825,II26824,WX8760);
	nand 	XG6668 	(II26794,II26793,WX8760);
	nand 	XG6669 	(II26763,II26762,WX8760);
	nand 	XG6670 	(II26732,II26731,WX8760);
	nand 	XG6671 	(II26701,II26700,WX8760);
	nand 	XG6672 	(II26670,II26669,WX8760);
	nand 	XG6673 	(II26639,II26638,WX8760);
	nand 	XG6674 	(II26608,II26607,WX8760);
	nand 	XG6675 	(II26577,II26576,WX8760);
	nand 	XG6676 	(II26546,II26545,WX8760);
	nand 	XG6677 	(II26515,II26514,WX8760);
	nand 	XG6678 	(II22975,II22974,WX7467);
	nand 	XG6679 	(II22944,II22943,WX7467);
	nand 	XG6680 	(II22913,II22912,WX7467);
	nand 	XG6681 	(II22882,II22881,WX7467);
	nand 	XG6682 	(II22851,II22850,WX7467);
	nand 	XG6683 	(II22820,II22819,WX7467);
	nand 	XG6684 	(II22789,II22788,WX7467);
	nand 	XG6685 	(II22758,II22757,WX7467);
	nand 	XG6686 	(II22727,II22726,WX7467);
	nand 	XG6687 	(II22696,II22695,WX7467);
	nand 	XG6688 	(II22665,II22664,WX7467);
	nand 	XG6689 	(II22634,II22633,WX7467);
	nand 	XG6690 	(II22603,II22602,WX7467);
	nand 	XG6691 	(II22572,II22571,WX7467);
	nand 	XG6692 	(II22541,II22540,WX7467);
	nand 	XG6693 	(II22510,II22509,WX7467);
	nand 	XG6694 	(II18970,II18969,WX6174);
	nand 	XG6695 	(II18939,II18938,WX6174);
	nand 	XG6696 	(II18908,II18907,WX6174);
	nand 	XG6697 	(II18877,II18876,WX6174);
	nand 	XG6698 	(II18846,II18845,WX6174);
	nand 	XG6699 	(II18815,II18814,WX6174);
	nand 	XG6700 	(II18784,II18783,WX6174);
	nand 	XG6701 	(II18753,II18752,WX6174);
	nand 	XG6702 	(II18722,II18721,WX6174);
	nand 	XG6703 	(II18691,II18690,WX6174);
	nand 	XG6704 	(II18660,II18659,WX6174);
	nand 	XG6705 	(II18629,II18628,WX6174);
	nand 	XG6706 	(II18598,II18597,WX6174);
	nand 	XG6707 	(II18567,II18566,WX6174);
	nand 	XG6708 	(II18536,II18535,WX6174);
	nand 	XG6709 	(II18505,II18504,WX6174);
	nand 	XG6710 	(II14965,II14964,WX4881);
	nand 	XG6711 	(II14934,II14933,WX4881);
	nand 	XG6712 	(II14903,II14902,WX4881);
	nand 	XG6713 	(II14872,II14871,WX4881);
	nand 	XG6714 	(II14841,II14840,WX4881);
	nand 	XG6715 	(II14810,II14809,WX4881);
	nand 	XG6716 	(II14779,II14778,WX4881);
	nand 	XG6717 	(II14748,II14747,WX4881);
	nand 	XG6718 	(II14717,II14716,WX4881);
	nand 	XG6719 	(II14686,II14685,WX4881);
	nand 	XG6720 	(II14655,II14654,WX4881);
	nand 	XG6721 	(II14624,II14623,WX4881);
	nand 	XG6722 	(II14593,II14592,WX4881);
	nand 	XG6723 	(II14562,II14561,WX4881);
	nand 	XG6724 	(II14531,II14530,WX4881);
	nand 	XG6725 	(II14500,II14499,WX4881);
	nand 	XG6726 	(II10960,II10959,WX3588);
	nand 	XG6727 	(II10929,II10928,WX3588);
	nand 	XG6728 	(II10898,II10897,WX3588);
	nand 	XG6729 	(II10867,II10866,WX3588);
	nand 	XG6730 	(II10836,II10835,WX3588);
	nand 	XG6731 	(II10805,II10804,WX3588);
	nand 	XG6732 	(II10774,II10773,WX3588);
	nand 	XG6733 	(II10743,II10742,WX3588);
	nand 	XG6734 	(II10712,II10711,WX3588);
	nand 	XG6735 	(II10681,II10680,WX3588);
	nand 	XG6736 	(II10650,II10649,WX3588);
	nand 	XG6737 	(II10619,II10618,WX3588);
	nand 	XG6738 	(II10588,II10587,WX3588);
	nand 	XG6739 	(II10557,II10556,WX3588);
	nand 	XG6740 	(II10526,II10525,WX3588);
	nand 	XG6741 	(II10495,II10494,WX3588);
	nand 	XG6742 	(II6955,II6954,WX2295);
	nand 	XG6743 	(II6924,II6923,WX2295);
	nand 	XG6744 	(II6893,II6892,WX2295);
	nand 	XG6745 	(II6862,II6861,WX2295);
	nand 	XG6746 	(II6831,II6830,WX2295);
	nand 	XG6747 	(II6800,II6799,WX2295);
	nand 	XG6748 	(II6769,II6768,WX2295);
	nand 	XG6749 	(II6738,II6737,WX2295);
	nand 	XG6750 	(II6707,II6706,WX2295);
	nand 	XG6751 	(II6676,II6675,WX2295);
	nand 	XG6752 	(II6645,II6644,WX2295);
	nand 	XG6753 	(II6614,II6613,WX2295);
	nand 	XG6754 	(II6583,II6582,WX2295);
	nand 	XG6755 	(II6552,II6551,WX2295);
	nand 	XG6756 	(II6521,II6520,WX2295);
	nand 	XG6757 	(II6490,II6489,WX2295);
	nand 	XG6758 	(II2950,II2949,WX1002);
	nand 	XG6759 	(II2919,II2918,WX1002);
	nand 	XG6760 	(II2888,II2887,WX1002);
	nand 	XG6761 	(II2857,II2856,WX1002);
	nand 	XG6762 	(II2826,II2825,WX1002);
	nand 	XG6763 	(II2795,II2794,WX1002);
	nand 	XG6764 	(II2764,II2763,WX1002);
	nand 	XG6765 	(II2733,II2732,WX1002);
	nand 	XG6766 	(II2702,II2701,WX1002);
	nand 	XG6767 	(II2671,II2670,WX1002);
	nand 	XG6768 	(II2640,II2639,WX1002);
	nand 	XG6769 	(II2609,II2608,WX1002);
	nand 	XG6770 	(II2578,II2577,WX1002);
	nand 	XG6771 	(II2547,II2546,WX1002);
	nand 	XG6772 	(II2516,II2515,WX1002);
	nand 	XG6773 	(II2485,II2484,WX1002);
	nand 	XG6774 	(II1990,II1988,WX645);
	nand 	XG6775 	(II2021,II2019,WX647);
	nand 	XG6776 	(II2052,II2050,WX649);
	nand 	XG6777 	(II2083,II2081,WX651);
	nand 	XG6778 	(II2114,II2112,WX653);
	nand 	XG6779 	(II2145,II2143,WX655);
	nand 	XG6780 	(II2176,II2174,WX657);
	nand 	XG6781 	(II2207,II2205,WX659);
	nand 	XG6782 	(II2238,II2236,WX661);
	nand 	XG6783 	(II2269,II2267,WX663);
	nand 	XG6784 	(II2300,II2298,WX665);
	nand 	XG6785 	(II2331,II2329,WX667);
	nand 	XG6786 	(II2362,II2360,WX669);
	nand 	XG6787 	(II2393,II2391,WX671);
	nand 	XG6788 	(II2424,II2422,WX673);
	nand 	XG6789 	(II2455,II2453,WX675);
	nand 	XG6790 	(II2486,II2484,WX677);
	nand 	XG6791 	(II2517,II2515,WX679);
	nand 	XG6792 	(II2548,II2546,WX681);
	nand 	XG6793 	(II2579,II2577,WX683);
	nand 	XG6794 	(II2610,II2608,WX685);
	nand 	XG6795 	(II2641,II2639,WX687);
	nand 	XG6796 	(II2672,II2670,WX689);
	nand 	XG6797 	(II2703,II2701,WX691);
	nand 	XG6798 	(II2734,II2732,WX693);
	nand 	XG6799 	(II2765,II2763,WX695);
	nand 	XG6800 	(II2796,II2794,WX697);
	nand 	XG6801 	(II2827,II2825,WX699);
	nand 	XG6802 	(II2858,II2856,WX701);
	nand 	XG6803 	(II2889,II2887,WX703);
	nand 	XG6804 	(II2920,II2918,WX705);
	nand 	XG6805 	(II2951,II2949,WX707);
	nand 	XG6806 	(II2002,II2005,II2004);
	nand 	XG6807 	(II2033,II2036,II2035);
	nand 	XG6808 	(II2064,II2067,II2066);
	nand 	XG6809 	(II2095,II2098,II2097);
	nand 	XG6810 	(II2126,II2129,II2128);
	nand 	XG6811 	(II2157,II2160,II2159);
	nand 	XG6812 	(II2188,II2191,II2190);
	nand 	XG6813 	(II2219,II2222,II2221);
	nand 	XG6814 	(II2250,II2253,II2252);
	nand 	XG6815 	(II2281,II2284,II2283);
	nand 	XG6816 	(II2312,II2315,II2314);
	nand 	XG6817 	(II2343,II2346,II2345);
	nand 	XG6818 	(II2374,II2377,II2376);
	nand 	XG6819 	(II2405,II2408,II2407);
	nand 	XG6820 	(II2436,II2439,II2438);
	nand 	XG6821 	(II2467,II2470,II2469);
	nand 	XG6822 	(II2498,II2501,II2500);
	nand 	XG6823 	(II2529,II2532,II2531);
	nand 	XG6824 	(II2560,II2563,II2562);
	nand 	XG6825 	(II2591,II2594,II2593);
	nand 	XG6826 	(II2622,II2625,II2624);
	nand 	XG6827 	(II2653,II2656,II2655);
	nand 	XG6828 	(II2684,II2687,II2686);
	nand 	XG6829 	(II2715,II2718,II2717);
	nand 	XG6830 	(II2746,II2749,II2748);
	nand 	XG6831 	(II2777,II2780,II2779);
	nand 	XG6832 	(II2808,II2811,II2810);
	nand 	XG6833 	(II2839,II2842,II2841);
	nand 	XG6834 	(II2870,II2873,II2872);
	nand 	XG6835 	(II2901,II2904,II2903);
	nand 	XG6836 	(II2932,II2935,II2934);
	nand 	XG6837 	(II2963,II2966,II2965);
	nand 	XG6838 	(II5995,II5993,WX1938);
	nand 	XG6839 	(II6026,II6024,WX1940);
	nand 	XG6840 	(II6057,II6055,WX1942);
	nand 	XG6841 	(II6088,II6086,WX1944);
	nand 	XG6842 	(II6119,II6117,WX1946);
	nand 	XG6843 	(II6150,II6148,WX1948);
	nand 	XG6844 	(II6181,II6179,WX1950);
	nand 	XG6845 	(II6212,II6210,WX1952);
	nand 	XG6846 	(II6243,II6241,WX1954);
	nand 	XG6847 	(II6274,II6272,WX1956);
	nand 	XG6848 	(II6305,II6303,WX1958);
	nand 	XG6849 	(II6336,II6334,WX1960);
	nand 	XG6850 	(II6367,II6365,WX1962);
	nand 	XG6851 	(II6398,II6396,WX1964);
	nand 	XG6852 	(II6429,II6427,WX1966);
	nand 	XG6853 	(II6460,II6458,WX1968);
	nand 	XG6854 	(II6491,II6489,WX1970);
	nand 	XG6855 	(II6522,II6520,WX1972);
	nand 	XG6856 	(II6553,II6551,WX1974);
	nand 	XG6857 	(II6584,II6582,WX1976);
	nand 	XG6858 	(II6615,II6613,WX1978);
	nand 	XG6859 	(II6646,II6644,WX1980);
	nand 	XG6860 	(II6677,II6675,WX1982);
	nand 	XG6861 	(II6708,II6706,WX1984);
	nand 	XG6862 	(II6739,II6737,WX1986);
	nand 	XG6863 	(II6770,II6768,WX1988);
	nand 	XG6864 	(II6801,II6799,WX1990);
	nand 	XG6865 	(II6832,II6830,WX1992);
	nand 	XG6866 	(II6863,II6861,WX1994);
	nand 	XG6867 	(II6894,II6892,WX1996);
	nand 	XG6868 	(II6925,II6923,WX1998);
	nand 	XG6869 	(II6956,II6954,WX2000);
	nand 	XG6870 	(II6007,II6010,II6009);
	nand 	XG6871 	(II6038,II6041,II6040);
	nand 	XG6872 	(II6069,II6072,II6071);
	nand 	XG6873 	(II6100,II6103,II6102);
	nand 	XG6874 	(II6131,II6134,II6133);
	nand 	XG6875 	(II6162,II6165,II6164);
	nand 	XG6876 	(II6193,II6196,II6195);
	nand 	XG6877 	(II6224,II6227,II6226);
	nand 	XG6878 	(II6255,II6258,II6257);
	nand 	XG6879 	(II6286,II6289,II6288);
	nand 	XG6880 	(II6317,II6320,II6319);
	nand 	XG6881 	(II6348,II6351,II6350);
	nand 	XG6882 	(II6379,II6382,II6381);
	nand 	XG6883 	(II6410,II6413,II6412);
	nand 	XG6884 	(II6441,II6444,II6443);
	nand 	XG6885 	(II6472,II6475,II6474);
	nand 	XG6886 	(II6503,II6506,II6505);
	nand 	XG6887 	(II6534,II6537,II6536);
	nand 	XG6888 	(II6565,II6568,II6567);
	nand 	XG6889 	(II6596,II6599,II6598);
	nand 	XG6890 	(II6627,II6630,II6629);
	nand 	XG6891 	(II6658,II6661,II6660);
	nand 	XG6892 	(II6689,II6692,II6691);
	nand 	XG6893 	(II6720,II6723,II6722);
	nand 	XG6894 	(II6751,II6754,II6753);
	nand 	XG6895 	(II6782,II6785,II6784);
	nand 	XG6896 	(II6813,II6816,II6815);
	nand 	XG6897 	(II6844,II6847,II6846);
	nand 	XG6898 	(II6875,II6878,II6877);
	nand 	XG6899 	(II6906,II6909,II6908);
	nand 	XG6900 	(II6937,II6940,II6939);
	nand 	XG6901 	(II6968,II6971,II6970);
	nand 	XG6902 	(II10000,II9998,WX3231);
	nand 	XG6903 	(II10031,II10029,WX3233);
	nand 	XG6904 	(II10062,II10060,WX3235);
	nand 	XG6905 	(II10093,II10091,WX3237);
	nand 	XG6906 	(II10124,II10122,WX3239);
	nand 	XG6907 	(II10155,II10153,WX3241);
	nand 	XG6908 	(II10186,II10184,WX3243);
	nand 	XG6909 	(II10217,II10215,WX3245);
	nand 	XG6910 	(II10248,II10246,WX3247);
	nand 	XG6911 	(II10279,II10277,WX3249);
	nand 	XG6912 	(II10310,II10308,WX3251);
	nand 	XG6913 	(II10341,II10339,WX3253);
	nand 	XG6914 	(II10372,II10370,WX3255);
	nand 	XG6915 	(II10403,II10401,WX3257);
	nand 	XG6916 	(II10434,II10432,WX3259);
	nand 	XG6917 	(II10465,II10463,WX3261);
	nand 	XG6918 	(II10496,II10494,WX3263);
	nand 	XG6919 	(II10527,II10525,WX3265);
	nand 	XG6920 	(II10558,II10556,WX3267);
	nand 	XG6921 	(II10589,II10587,WX3269);
	nand 	XG6922 	(II10620,II10618,WX3271);
	nand 	XG6923 	(II10651,II10649,WX3273);
	nand 	XG6924 	(II10682,II10680,WX3275);
	nand 	XG6925 	(II10713,II10711,WX3277);
	nand 	XG6926 	(II10744,II10742,WX3279);
	nand 	XG6927 	(II10775,II10773,WX3281);
	nand 	XG6928 	(II10806,II10804,WX3283);
	nand 	XG6929 	(II10837,II10835,WX3285);
	nand 	XG6930 	(II10868,II10866,WX3287);
	nand 	XG6931 	(II10899,II10897,WX3289);
	nand 	XG6932 	(II10930,II10928,WX3291);
	nand 	XG6933 	(II10961,II10959,WX3293);
	nand 	XG6934 	(II10012,II10015,II10014);
	nand 	XG6935 	(II10043,II10046,II10045);
	nand 	XG6936 	(II10074,II10077,II10076);
	nand 	XG6937 	(II10105,II10108,II10107);
	nand 	XG6938 	(II10136,II10139,II10138);
	nand 	XG6939 	(II10167,II10170,II10169);
	nand 	XG6940 	(II10198,II10201,II10200);
	nand 	XG6941 	(II10229,II10232,II10231);
	nand 	XG6942 	(II10260,II10263,II10262);
	nand 	XG6943 	(II10291,II10294,II10293);
	nand 	XG6944 	(II10322,II10325,II10324);
	nand 	XG6945 	(II10353,II10356,II10355);
	nand 	XG6946 	(II10384,II10387,II10386);
	nand 	XG6947 	(II10415,II10418,II10417);
	nand 	XG6948 	(II10446,II10449,II10448);
	nand 	XG6949 	(II10477,II10480,II10479);
	nand 	XG6950 	(II10508,II10511,II10510);
	nand 	XG6951 	(II10539,II10542,II10541);
	nand 	XG6952 	(II10570,II10573,II10572);
	nand 	XG6953 	(II10601,II10604,II10603);
	nand 	XG6954 	(II10632,II10635,II10634);
	nand 	XG6955 	(II10663,II10666,II10665);
	nand 	XG6956 	(II10694,II10697,II10696);
	nand 	XG6957 	(II10725,II10728,II10727);
	nand 	XG6958 	(II10756,II10759,II10758);
	nand 	XG6959 	(II10787,II10790,II10789);
	nand 	XG6960 	(II10818,II10821,II10820);
	nand 	XG6961 	(II10849,II10852,II10851);
	nand 	XG6962 	(II10880,II10883,II10882);
	nand 	XG6963 	(II10911,II10914,II10913);
	nand 	XG6964 	(II10942,II10945,II10944);
	nand 	XG6965 	(II10973,II10976,II10975);
	nand 	XG6966 	(II14005,II14003,WX4524);
	nand 	XG6967 	(II14036,II14034,WX4526);
	nand 	XG6968 	(II14067,II14065,WX4528);
	nand 	XG6969 	(II14098,II14096,WX4530);
	nand 	XG6970 	(II14129,II14127,WX4532);
	nand 	XG6971 	(II14160,II14158,WX4534);
	nand 	XG6972 	(II14191,II14189,WX4536);
	nand 	XG6973 	(II14222,II14220,WX4538);
	nand 	XG6974 	(II14253,II14251,WX4540);
	nand 	XG6975 	(II14284,II14282,WX4542);
	nand 	XG6976 	(II14315,II14313,WX4544);
	nand 	XG6977 	(II14346,II14344,WX4546);
	nand 	XG6978 	(II14377,II14375,WX4548);
	nand 	XG6979 	(II14408,II14406,WX4550);
	nand 	XG6980 	(II14439,II14437,WX4552);
	nand 	XG6981 	(II14470,II14468,WX4554);
	nand 	XG6982 	(II14501,II14499,WX4556);
	nand 	XG6983 	(II14532,II14530,WX4558);
	nand 	XG6984 	(II14563,II14561,WX4560);
	nand 	XG6985 	(II14594,II14592,WX4562);
	nand 	XG6986 	(II14625,II14623,WX4564);
	nand 	XG6987 	(II14656,II14654,WX4566);
	nand 	XG6988 	(II14687,II14685,WX4568);
	nand 	XG6989 	(II14718,II14716,WX4570);
	nand 	XG6990 	(II14749,II14747,WX4572);
	nand 	XG6991 	(II14780,II14778,WX4574);
	nand 	XG6992 	(II14811,II14809,WX4576);
	nand 	XG6993 	(II14842,II14840,WX4578);
	nand 	XG6994 	(II14873,II14871,WX4580);
	nand 	XG6995 	(II14904,II14902,WX4582);
	nand 	XG6996 	(II14935,II14933,WX4584);
	nand 	XG6997 	(II14966,II14964,WX4586);
	nand 	XG6998 	(II14017,II14020,II14019);
	nand 	XG6999 	(II14048,II14051,II14050);
	nand 	XG7000 	(II14079,II14082,II14081);
	nand 	XG7001 	(II14110,II14113,II14112);
	nand 	XG7002 	(II14141,II14144,II14143);
	nand 	XG7003 	(II14172,II14175,II14174);
	nand 	XG7004 	(II14203,II14206,II14205);
	nand 	XG7005 	(II14234,II14237,II14236);
	nand 	XG7006 	(II14265,II14268,II14267);
	nand 	XG7007 	(II14296,II14299,II14298);
	nand 	XG7008 	(II14327,II14330,II14329);
	nand 	XG7009 	(II14358,II14361,II14360);
	nand 	XG7010 	(II14389,II14392,II14391);
	nand 	XG7011 	(II14420,II14423,II14422);
	nand 	XG7012 	(II14451,II14454,II14453);
	nand 	XG7013 	(II14482,II14485,II14484);
	nand 	XG7014 	(II14513,II14516,II14515);
	nand 	XG7015 	(II14544,II14547,II14546);
	nand 	XG7016 	(II14575,II14578,II14577);
	nand 	XG7017 	(II14606,II14609,II14608);
	nand 	XG7018 	(II14637,II14640,II14639);
	nand 	XG7019 	(II14668,II14671,II14670);
	nand 	XG7020 	(II14699,II14702,II14701);
	nand 	XG7021 	(II14730,II14733,II14732);
	nand 	XG7022 	(II14761,II14764,II14763);
	nand 	XG7023 	(II14792,II14795,II14794);
	nand 	XG7024 	(II14823,II14826,II14825);
	nand 	XG7025 	(II14854,II14857,II14856);
	nand 	XG7026 	(II14885,II14888,II14887);
	nand 	XG7027 	(II14916,II14919,II14918);
	nand 	XG7028 	(II14947,II14950,II14949);
	nand 	XG7029 	(II14978,II14981,II14980);
	nand 	XG7030 	(II18010,II18008,WX5817);
	nand 	XG7031 	(II18041,II18039,WX5819);
	nand 	XG7032 	(II18072,II18070,WX5821);
	nand 	XG7033 	(II18103,II18101,WX5823);
	nand 	XG7034 	(II18134,II18132,WX5825);
	nand 	XG7035 	(II18165,II18163,WX5827);
	nand 	XG7036 	(II18196,II18194,WX5829);
	nand 	XG7037 	(II18227,II18225,WX5831);
	nand 	XG7038 	(II18258,II18256,WX5833);
	nand 	XG7039 	(II18289,II18287,WX5835);
	nand 	XG7040 	(II18320,II18318,WX5837);
	nand 	XG7041 	(II18351,II18349,WX5839);
	nand 	XG7042 	(II18382,II18380,WX5841);
	nand 	XG7043 	(II18413,II18411,WX5843);
	nand 	XG7044 	(II18444,II18442,WX5845);
	nand 	XG7045 	(II18475,II18473,WX5847);
	nand 	XG7046 	(II18506,II18504,WX5849);
	nand 	XG7047 	(II18537,II18535,WX5851);
	nand 	XG7048 	(II18568,II18566,WX5853);
	nand 	XG7049 	(II18599,II18597,WX5855);
	nand 	XG7050 	(II18630,II18628,WX5857);
	nand 	XG7051 	(II18661,II18659,WX5859);
	nand 	XG7052 	(II18692,II18690,WX5861);
	nand 	XG7053 	(II18723,II18721,WX5863);
	nand 	XG7054 	(II18754,II18752,WX5865);
	nand 	XG7055 	(II18785,II18783,WX5867);
	nand 	XG7056 	(II18816,II18814,WX5869);
	nand 	XG7057 	(II18847,II18845,WX5871);
	nand 	XG7058 	(II18878,II18876,WX5873);
	nand 	XG7059 	(II18909,II18907,WX5875);
	nand 	XG7060 	(II18940,II18938,WX5877);
	nand 	XG7061 	(II18971,II18969,WX5879);
	nand 	XG7062 	(II18022,II18025,II18024);
	nand 	XG7063 	(II18053,II18056,II18055);
	nand 	XG7064 	(II18084,II18087,II18086);
	nand 	XG7065 	(II18115,II18118,II18117);
	nand 	XG7066 	(II18146,II18149,II18148);
	nand 	XG7067 	(II18177,II18180,II18179);
	nand 	XG7068 	(II18208,II18211,II18210);
	nand 	XG7069 	(II18239,II18242,II18241);
	nand 	XG7070 	(II18270,II18273,II18272);
	nand 	XG7071 	(II18301,II18304,II18303);
	nand 	XG7072 	(II18332,II18335,II18334);
	nand 	XG7073 	(II18363,II18366,II18365);
	nand 	XG7074 	(II18394,II18397,II18396);
	nand 	XG7075 	(II18425,II18428,II18427);
	nand 	XG7076 	(II18456,II18459,II18458);
	nand 	XG7077 	(II18487,II18490,II18489);
	nand 	XG7078 	(II18518,II18521,II18520);
	nand 	XG7079 	(II18549,II18552,II18551);
	nand 	XG7080 	(II18580,II18583,II18582);
	nand 	XG7081 	(II18611,II18614,II18613);
	nand 	XG7082 	(II18642,II18645,II18644);
	nand 	XG7083 	(II18673,II18676,II18675);
	nand 	XG7084 	(II18704,II18707,II18706);
	nand 	XG7085 	(II18735,II18738,II18737);
	nand 	XG7086 	(II18766,II18769,II18768);
	nand 	XG7087 	(II18797,II18800,II18799);
	nand 	XG7088 	(II18828,II18831,II18830);
	nand 	XG7089 	(II18859,II18862,II18861);
	nand 	XG7090 	(II18890,II18893,II18892);
	nand 	XG7091 	(II18921,II18924,II18923);
	nand 	XG7092 	(II18952,II18955,II18954);
	nand 	XG7093 	(II18983,II18986,II18985);
	nand 	XG7094 	(II22015,II22013,WX7110);
	nand 	XG7095 	(II22046,II22044,WX7112);
	nand 	XG7096 	(II22077,II22075,WX7114);
	nand 	XG7097 	(II22108,II22106,WX7116);
	nand 	XG7098 	(II22139,II22137,WX7118);
	nand 	XG7099 	(II22170,II22168,WX7120);
	nand 	XG7100 	(II22201,II22199,WX7122);
	nand 	XG7101 	(II22232,II22230,WX7124);
	nand 	XG7102 	(II22263,II22261,WX7126);
	nand 	XG7103 	(II22294,II22292,WX7128);
	nand 	XG7104 	(II22325,II22323,WX7130);
	nand 	XG7105 	(II22356,II22354,WX7132);
	nand 	XG7106 	(II22387,II22385,WX7134);
	nand 	XG7107 	(II22418,II22416,WX7136);
	nand 	XG7108 	(II22449,II22447,WX7138);
	nand 	XG7109 	(II22480,II22478,WX7140);
	nand 	XG7110 	(II22511,II22509,WX7142);
	nand 	XG7111 	(II22542,II22540,WX7144);
	nand 	XG7112 	(II22573,II22571,WX7146);
	nand 	XG7113 	(II22604,II22602,WX7148);
	nand 	XG7114 	(II22635,II22633,WX7150);
	nand 	XG7115 	(II22666,II22664,WX7152);
	nand 	XG7116 	(II22697,II22695,WX7154);
	nand 	XG7117 	(II22728,II22726,WX7156);
	nand 	XG7118 	(II22759,II22757,WX7158);
	nand 	XG7119 	(II22790,II22788,WX7160);
	nand 	XG7120 	(II22821,II22819,WX7162);
	nand 	XG7121 	(II22852,II22850,WX7164);
	nand 	XG7122 	(II22883,II22881,WX7166);
	nand 	XG7123 	(II22914,II22912,WX7168);
	nand 	XG7124 	(II22945,II22943,WX7170);
	nand 	XG7125 	(II22976,II22974,WX7172);
	nand 	XG7126 	(II22027,II22030,II22029);
	nand 	XG7127 	(II22058,II22061,II22060);
	nand 	XG7128 	(II22089,II22092,II22091);
	nand 	XG7129 	(II22120,II22123,II22122);
	nand 	XG7130 	(II22151,II22154,II22153);
	nand 	XG7131 	(II22182,II22185,II22184);
	nand 	XG7132 	(II22213,II22216,II22215);
	nand 	XG7133 	(II22244,II22247,II22246);
	nand 	XG7134 	(II22275,II22278,II22277);
	nand 	XG7135 	(II22306,II22309,II22308);
	nand 	XG7136 	(II22337,II22340,II22339);
	nand 	XG7137 	(II22368,II22371,II22370);
	nand 	XG7138 	(II22399,II22402,II22401);
	nand 	XG7139 	(II22430,II22433,II22432);
	nand 	XG7140 	(II22461,II22464,II22463);
	nand 	XG7141 	(II22492,II22495,II22494);
	nand 	XG7142 	(II22523,II22526,II22525);
	nand 	XG7143 	(II22554,II22557,II22556);
	nand 	XG7144 	(II22585,II22588,II22587);
	nand 	XG7145 	(II22616,II22619,II22618);
	nand 	XG7146 	(II22647,II22650,II22649);
	nand 	XG7147 	(II22678,II22681,II22680);
	nand 	XG7148 	(II22709,II22712,II22711);
	nand 	XG7149 	(II22740,II22743,II22742);
	nand 	XG7150 	(II22771,II22774,II22773);
	nand 	XG7151 	(II22802,II22805,II22804);
	nand 	XG7152 	(II22833,II22836,II22835);
	nand 	XG7153 	(II22864,II22867,II22866);
	nand 	XG7154 	(II22895,II22898,II22897);
	nand 	XG7155 	(II22926,II22929,II22928);
	nand 	XG7156 	(II22957,II22960,II22959);
	nand 	XG7157 	(II22988,II22991,II22990);
	nand 	XG7158 	(II26020,II26018,WX8403);
	nand 	XG7159 	(II26051,II26049,WX8405);
	nand 	XG7160 	(II26082,II26080,WX8407);
	nand 	XG7161 	(II26113,II26111,WX8409);
	nand 	XG7162 	(II26144,II26142,WX8411);
	nand 	XG7163 	(II26175,II26173,WX8413);
	nand 	XG7164 	(II26206,II26204,WX8415);
	nand 	XG7165 	(II26237,II26235,WX8417);
	nand 	XG7166 	(II26268,II26266,WX8419);
	nand 	XG7167 	(II26299,II26297,WX8421);
	nand 	XG7168 	(II26330,II26328,WX8423);
	nand 	XG7169 	(II26361,II26359,WX8425);
	nand 	XG7170 	(II26392,II26390,WX8427);
	nand 	XG7171 	(II26423,II26421,WX8429);
	nand 	XG7172 	(II26454,II26452,WX8431);
	nand 	XG7173 	(II26485,II26483,WX8433);
	nand 	XG7174 	(II26516,II26514,WX8435);
	nand 	XG7175 	(II26547,II26545,WX8437);
	nand 	XG7176 	(II26578,II26576,WX8439);
	nand 	XG7177 	(II26609,II26607,WX8441);
	nand 	XG7178 	(II26640,II26638,WX8443);
	nand 	XG7179 	(II26671,II26669,WX8445);
	nand 	XG7180 	(II26702,II26700,WX8447);
	nand 	XG7181 	(II26733,II26731,WX8449);
	nand 	XG7182 	(II26764,II26762,WX8451);
	nand 	XG7183 	(II26795,II26793,WX8453);
	nand 	XG7184 	(II26826,II26824,WX8455);
	nand 	XG7185 	(II26857,II26855,WX8457);
	nand 	XG7186 	(II26888,II26886,WX8459);
	nand 	XG7187 	(II26919,II26917,WX8461);
	nand 	XG7188 	(II26950,II26948,WX8463);
	nand 	XG7189 	(II26981,II26979,WX8465);
	nand 	XG7190 	(II26032,II26035,II26034);
	nand 	XG7191 	(II26063,II26066,II26065);
	nand 	XG7192 	(II26094,II26097,II26096);
	nand 	XG7193 	(II26125,II26128,II26127);
	nand 	XG7194 	(II26156,II26159,II26158);
	nand 	XG7195 	(II26187,II26190,II26189);
	nand 	XG7196 	(II26218,II26221,II26220);
	nand 	XG7197 	(II26249,II26252,II26251);
	nand 	XG7198 	(II26280,II26283,II26282);
	nand 	XG7199 	(II26311,II26314,II26313);
	nand 	XG7200 	(II26342,II26345,II26344);
	nand 	XG7201 	(II26373,II26376,II26375);
	nand 	XG7202 	(II26404,II26407,II26406);
	nand 	XG7203 	(II26435,II26438,II26437);
	nand 	XG7204 	(II26466,II26469,II26468);
	nand 	XG7205 	(II26497,II26500,II26499);
	nand 	XG7206 	(II26528,II26531,II26530);
	nand 	XG7207 	(II26559,II26562,II26561);
	nand 	XG7208 	(II26590,II26593,II26592);
	nand 	XG7209 	(II26621,II26624,II26623);
	nand 	XG7210 	(II26652,II26655,II26654);
	nand 	XG7211 	(II26683,II26686,II26685);
	nand 	XG7212 	(II26714,II26717,II26716);
	nand 	XG7213 	(II26745,II26748,II26747);
	nand 	XG7214 	(II26776,II26779,II26778);
	nand 	XG7215 	(II26807,II26810,II26809);
	nand 	XG7216 	(II26838,II26841,II26840);
	nand 	XG7217 	(II26869,II26872,II26871);
	nand 	XG7218 	(II26900,II26903,II26902);
	nand 	XG7219 	(II26931,II26934,II26933);
	nand 	XG7220 	(II26962,II26965,II26964);
	nand 	XG7221 	(II26993,II26996,II26995);
	nand 	XG7222 	(II30025,II30023,WX9696);
	nand 	XG7223 	(II30056,II30054,WX9698);
	nand 	XG7224 	(II30087,II30085,WX9700);
	nand 	XG7225 	(II30118,II30116,WX9702);
	nand 	XG7226 	(II30149,II30147,WX9704);
	nand 	XG7227 	(II30180,II30178,WX9706);
	nand 	XG7228 	(II30211,II30209,WX9708);
	nand 	XG7229 	(II30242,II30240,WX9710);
	nand 	XG7230 	(II30273,II30271,WX9712);
	nand 	XG7231 	(II30304,II30302,WX9714);
	nand 	XG7232 	(II30335,II30333,WX9716);
	nand 	XG7233 	(II30366,II30364,WX9718);
	nand 	XG7234 	(II30397,II30395,WX9720);
	nand 	XG7235 	(II30428,II30426,WX9722);
	nand 	XG7236 	(II30459,II30457,WX9724);
	nand 	XG7237 	(II30490,II30488,WX9726);
	nand 	XG7238 	(II30521,II30519,WX9728);
	nand 	XG7239 	(II30552,II30550,WX9730);
	nand 	XG7240 	(II30583,II30581,WX9732);
	nand 	XG7241 	(II30614,II30612,WX9734);
	nand 	XG7242 	(II30645,II30643,WX9736);
	nand 	XG7243 	(II30676,II30674,WX9738);
	nand 	XG7244 	(II30707,II30705,WX9740);
	nand 	XG7245 	(II30738,II30736,WX9742);
	nand 	XG7246 	(II30769,II30767,WX9744);
	nand 	XG7247 	(II30800,II30798,WX9746);
	nand 	XG7248 	(II30831,II30829,WX9748);
	nand 	XG7249 	(II30862,II30860,WX9750);
	nand 	XG7250 	(II30893,II30891,WX9752);
	nand 	XG7251 	(II30924,II30922,WX9754);
	nand 	XG7252 	(II30955,II30953,WX9756);
	nand 	XG7253 	(II30986,II30984,WX9758);
	nand 	XG7254 	(II30037,II30040,II30039);
	nand 	XG7255 	(II30068,II30071,II30070);
	nand 	XG7256 	(II30099,II30102,II30101);
	nand 	XG7257 	(II30130,II30133,II30132);
	nand 	XG7258 	(II30161,II30164,II30163);
	nand 	XG7259 	(II30192,II30195,II30194);
	nand 	XG7260 	(II30223,II30226,II30225);
	nand 	XG7261 	(II30254,II30257,II30256);
	nand 	XG7262 	(II30285,II30288,II30287);
	nand 	XG7263 	(II30316,II30319,II30318);
	nand 	XG7264 	(II30347,II30350,II30349);
	nand 	XG7265 	(II30378,II30381,II30380);
	nand 	XG7266 	(II30409,II30412,II30411);
	nand 	XG7267 	(II30440,II30443,II30442);
	nand 	XG7268 	(II30471,II30474,II30473);
	nand 	XG7269 	(II30502,II30505,II30504);
	nand 	XG7270 	(II30533,II30536,II30535);
	nand 	XG7271 	(II30564,II30567,II30566);
	nand 	XG7272 	(II30595,II30598,II30597);
	nand 	XG7273 	(II30626,II30629,II30628);
	nand 	XG7274 	(II30657,II30660,II30659);
	nand 	XG7275 	(II30688,II30691,II30690);
	nand 	XG7276 	(II30719,II30722,II30721);
	nand 	XG7277 	(II30750,II30753,II30752);
	nand 	XG7278 	(II30781,II30784,II30783);
	nand 	XG7279 	(II30812,II30815,II30814);
	nand 	XG7280 	(II30843,II30846,II30845);
	nand 	XG7281 	(II30874,II30877,II30876);
	nand 	XG7282 	(II30905,II30908,II30907);
	nand 	XG7283 	(II30936,II30939,II30938);
	nand 	XG7284 	(II30967,II30970,II30969);
	nand 	XG7285 	(II30998,II31001,II31000);
	nand 	XG7286 	(II34030,II34028,WX10989);
	nand 	XG7287 	(II34061,II34059,WX10991);
	nand 	XG7288 	(II34092,II34090,WX10993);
	nand 	XG7289 	(II34123,II34121,WX10995);
	nand 	XG7290 	(II34154,II34152,WX10997);
	nand 	XG7291 	(II34185,II34183,WX10999);
	nand 	XG7292 	(II34216,II34214,WX11001);
	nand 	XG7293 	(II34247,II34245,WX11003);
	nand 	XG7294 	(II34278,II34276,WX11005);
	nand 	XG7295 	(II34309,II34307,WX11007);
	nand 	XG7296 	(II34340,II34338,WX11009);
	nand 	XG7297 	(II34371,II34369,WX11011);
	nand 	XG7298 	(II34402,II34400,WX11013);
	nand 	XG7299 	(II34433,II34431,WX11015);
	nand 	XG7300 	(II34464,II34462,WX11017);
	nand 	XG7301 	(II34495,II34493,WX11019);
	nand 	XG7302 	(II34526,II34524,WX11021);
	nand 	XG7303 	(II34557,II34555,WX11023);
	nand 	XG7304 	(II34588,II34586,WX11025);
	nand 	XG7305 	(II34619,II34617,WX11027);
	nand 	XG7306 	(II34650,II34648,WX11029);
	nand 	XG7307 	(II34681,II34679,WX11031);
	nand 	XG7308 	(II34712,II34710,WX11033);
	nand 	XG7309 	(II34743,II34741,WX11035);
	nand 	XG7310 	(II34774,II34772,WX11037);
	nand 	XG7311 	(II34805,II34803,WX11039);
	nand 	XG7312 	(II34836,II34834,WX11041);
	nand 	XG7313 	(II34867,II34865,WX11043);
	nand 	XG7314 	(II34898,II34896,WX11045);
	nand 	XG7315 	(II34929,II34927,WX11047);
	nand 	XG7316 	(II34960,II34958,WX11049);
	nand 	XG7317 	(II34991,II34989,WX11051);
	nand 	XG7318 	(II34042,II34045,II34044);
	nand 	XG7319 	(II34073,II34076,II34075);
	nand 	XG7320 	(II34104,II34107,II34106);
	nand 	XG7321 	(II34135,II34138,II34137);
	nand 	XG7322 	(II34166,II34169,II34168);
	nand 	XG7323 	(II34197,II34200,II34199);
	nand 	XG7324 	(II34228,II34231,II34230);
	nand 	XG7325 	(II34259,II34262,II34261);
	nand 	XG7326 	(II34290,II34293,II34292);
	nand 	XG7327 	(II34321,II34324,II34323);
	nand 	XG7328 	(II34352,II34355,II34354);
	nand 	XG7329 	(II34383,II34386,II34385);
	nand 	XG7330 	(II34414,II34417,II34416);
	nand 	XG7331 	(II34445,II34448,II34447);
	nand 	XG7332 	(II34476,II34479,II34478);
	nand 	XG7333 	(II34507,II34510,II34509);
	nand 	XG7334 	(II34538,II34541,II34540);
	nand 	XG7335 	(II34569,II34572,II34571);
	nand 	XG7336 	(II34600,II34603,II34602);
	nand 	XG7337 	(II34631,II34634,II34633);
	nand 	XG7338 	(II34662,II34665,II34664);
	nand 	XG7339 	(II34693,II34696,II34695);
	nand 	XG7340 	(II34724,II34727,II34726);
	nand 	XG7341 	(II34755,II34758,II34757);
	nand 	XG7342 	(II34786,II34789,II34788);
	nand 	XG7343 	(II34817,II34820,II34819);
	nand 	XG7344 	(II34848,II34851,II34850);
	nand 	XG7345 	(II34879,II34882,II34881);
	nand 	XG7346 	(II34910,II34913,II34912);
	nand 	XG7347 	(II34941,II34944,II34943);
	nand 	XG7348 	(II34972,II34975,II34974);
	nand 	XG7349 	(II35003,II35006,II35005);
	nand 	XG7350 	(II35555,II35554,WX10987);
	nand 	XG7351 	(II35751,II35750,WX10986);
	nand 	XG7352 	(II35744,II35743,WX10985);
	nand 	XG7353 	(II35737,II35736,WX10984);
	nand 	XG7354 	(II35541,II35540,WX10983);
	nand 	XG7355 	(II35730,II35729,WX10982);
	nand 	XG7356 	(II35723,II35722,WX10981);
	nand 	XG7357 	(II35716,II35715,WX10980);
	nand 	XG7358 	(II35709,II35708,WX10979);
	nand 	XG7359 	(II35702,II35701,WX10978);
	nand 	XG7360 	(II35695,II35694,WX10977);
	nand 	XG7361 	(II35526,II35525,WX10976);
	nand 	XG7362 	(II35688,II35687,WX10975);
	nand 	XG7363 	(II35681,II35680,WX10974);
	nand 	XG7364 	(II35674,II35673,WX10973);
	nand 	XG7365 	(II35667,II35666,WX10972);
	nand 	XG7366 	(II35511,II35510,WX10971);
	nand 	XG7367 	(II35660,II35659,WX10970);
	nand 	XG7368 	(II35653,II35652,WX10969);
	nand 	XG7369 	(II35646,II35645,WX10968);
	nand 	XG7370 	(II35639,II35638,WX10967);
	nand 	XG7371 	(II35632,II35631,WX10966);
	nand 	XG7372 	(II35625,II35624,WX10965);
	nand 	XG7373 	(II35618,II35617,WX10964);
	nand 	XG7374 	(II35611,II35610,WX10963);
	nand 	XG7375 	(II35604,II35603,WX10962);
	nand 	XG7376 	(II35597,II35596,WX10961);
	nand 	XG7377 	(II35590,II35589,WX10960);
	nand 	XG7378 	(II35583,II35582,WX10959);
	nand 	XG7379 	(II35576,II35575,WX10958);
	nand 	XG7380 	(II35569,II35568,WX10957);
	nand 	XG7381 	(II35562,II35561,WX10956);
	nand 	XG7382 	(II31550,II31549,WX9694);
	nand 	XG7383 	(II31746,II31745,WX9693);
	nand 	XG7384 	(II31739,II31738,WX9692);
	nand 	XG7385 	(II31732,II31731,WX9691);
	nand 	XG7386 	(II31536,II31535,WX9690);
	nand 	XG7387 	(II31725,II31724,WX9689);
	nand 	XG7388 	(II31718,II31717,WX9688);
	nand 	XG7389 	(II31711,II31710,WX9687);
	nand 	XG7390 	(II31704,II31703,WX9686);
	nand 	XG7391 	(II31697,II31696,WX9685);
	nand 	XG7392 	(II31690,II31689,WX9684);
	nand 	XG7393 	(II31521,II31520,WX9683);
	nand 	XG7394 	(II31683,II31682,WX9682);
	nand 	XG7395 	(II31676,II31675,WX9681);
	nand 	XG7396 	(II31669,II31668,WX9680);
	nand 	XG7397 	(II31662,II31661,WX9679);
	nand 	XG7398 	(II31506,II31505,WX9678);
	nand 	XG7399 	(II31655,II31654,WX9677);
	nand 	XG7400 	(II31648,II31647,WX9676);
	nand 	XG7401 	(II31641,II31640,WX9675);
	nand 	XG7402 	(II31634,II31633,WX9674);
	nand 	XG7403 	(II31627,II31626,WX9673);
	nand 	XG7404 	(II31620,II31619,WX9672);
	nand 	XG7405 	(II31613,II31612,WX9671);
	nand 	XG7406 	(II31606,II31605,WX9670);
	nand 	XG7407 	(II31599,II31598,WX9669);
	nand 	XG7408 	(II31592,II31591,WX9668);
	nand 	XG7409 	(II31585,II31584,WX9667);
	nand 	XG7410 	(II31578,II31577,WX9666);
	nand 	XG7411 	(II31571,II31570,WX9665);
	nand 	XG7412 	(II31564,II31563,WX9664);
	nand 	XG7413 	(II31557,II31556,WX9663);
	nand 	XG7414 	(II27545,II27544,WX8401);
	nand 	XG7415 	(II27741,II27740,WX8400);
	nand 	XG7416 	(II27734,II27733,WX8399);
	nand 	XG7417 	(II27727,II27726,WX8398);
	nand 	XG7418 	(II27531,II27530,WX8397);
	nand 	XG7419 	(II27720,II27719,WX8396);
	nand 	XG7420 	(II27713,II27712,WX8395);
	nand 	XG7421 	(II27706,II27705,WX8394);
	nand 	XG7422 	(II27699,II27698,WX8393);
	nand 	XG7423 	(II27692,II27691,WX8392);
	nand 	XG7424 	(II27685,II27684,WX8391);
	nand 	XG7425 	(II27516,II27515,WX8390);
	nand 	XG7426 	(II27678,II27677,WX8389);
	nand 	XG7427 	(II27671,II27670,WX8388);
	nand 	XG7428 	(II27664,II27663,WX8387);
	nand 	XG7429 	(II27657,II27656,WX8386);
	nand 	XG7430 	(II27501,II27500,WX8385);
	nand 	XG7431 	(II27650,II27649,WX8384);
	nand 	XG7432 	(II27643,II27642,WX8383);
	nand 	XG7433 	(II27636,II27635,WX8382);
	nand 	XG7434 	(II27629,II27628,WX8381);
	nand 	XG7435 	(II27622,II27621,WX8380);
	nand 	XG7436 	(II27615,II27614,WX8379);
	nand 	XG7437 	(II27608,II27607,WX8378);
	nand 	XG7438 	(II27601,II27600,WX8377);
	nand 	XG7439 	(II27594,II27593,WX8376);
	nand 	XG7440 	(II27587,II27586,WX8375);
	nand 	XG7441 	(II27580,II27579,WX8374);
	nand 	XG7442 	(II27573,II27572,WX8373);
	nand 	XG7443 	(II27566,II27565,WX8372);
	nand 	XG7444 	(II27559,II27558,WX8371);
	nand 	XG7445 	(II27552,II27551,WX8370);
	nand 	XG7446 	(II23540,II23539,WX7108);
	nand 	XG7447 	(II23736,II23735,WX7107);
	nand 	XG7448 	(II23729,II23728,WX7106);
	nand 	XG7449 	(II23722,II23721,WX7105);
	nand 	XG7450 	(II23526,II23525,WX7104);
	nand 	XG7451 	(II23715,II23714,WX7103);
	nand 	XG7452 	(II23708,II23707,WX7102);
	nand 	XG7453 	(II23701,II23700,WX7101);
	nand 	XG7454 	(II23694,II23693,WX7100);
	nand 	XG7455 	(II23687,II23686,WX7099);
	nand 	XG7456 	(II23680,II23679,WX7098);
	nand 	XG7457 	(II23511,II23510,WX7097);
	nand 	XG7458 	(II23673,II23672,WX7096);
	nand 	XG7459 	(II23666,II23665,WX7095);
	nand 	XG7460 	(II23659,II23658,WX7094);
	nand 	XG7461 	(II23652,II23651,WX7093);
	nand 	XG7462 	(II23496,II23495,WX7092);
	nand 	XG7463 	(II23645,II23644,WX7091);
	nand 	XG7464 	(II23638,II23637,WX7090);
	nand 	XG7465 	(II23631,II23630,WX7089);
	nand 	XG7466 	(II23624,II23623,WX7088);
	nand 	XG7467 	(II23617,II23616,WX7087);
	nand 	XG7468 	(II23610,II23609,WX7086);
	nand 	XG7469 	(II23603,II23602,WX7085);
	nand 	XG7470 	(II23596,II23595,WX7084);
	nand 	XG7471 	(II23589,II23588,WX7083);
	nand 	XG7472 	(II23582,II23581,WX7082);
	nand 	XG7473 	(II23575,II23574,WX7081);
	nand 	XG7474 	(II23568,II23567,WX7080);
	nand 	XG7475 	(II23561,II23560,WX7079);
	nand 	XG7476 	(II23554,II23553,WX7078);
	nand 	XG7477 	(II23547,II23546,WX7077);
	nand 	XG7478 	(II19535,II19534,WX5815);
	nand 	XG7479 	(II19731,II19730,WX5814);
	nand 	XG7480 	(II19724,II19723,WX5813);
	nand 	XG7481 	(II19717,II19716,WX5812);
	nand 	XG7482 	(II19521,II19520,WX5811);
	nand 	XG7483 	(II19710,II19709,WX5810);
	nand 	XG7484 	(II19703,II19702,WX5809);
	nand 	XG7485 	(II19696,II19695,WX5808);
	nand 	XG7486 	(II19689,II19688,WX5807);
	nand 	XG7487 	(II19682,II19681,WX5806);
	nand 	XG7488 	(II19675,II19674,WX5805);
	nand 	XG7489 	(II19506,II19505,WX5804);
	nand 	XG7490 	(II19668,II19667,WX5803);
	nand 	XG7491 	(II19661,II19660,WX5802);
	nand 	XG7492 	(II19654,II19653,WX5801);
	nand 	XG7493 	(II19647,II19646,WX5800);
	nand 	XG7494 	(II19491,II19490,WX5799);
	nand 	XG7495 	(II19640,II19639,WX5798);
	nand 	XG7496 	(II19633,II19632,WX5797);
	nand 	XG7497 	(II19626,II19625,WX5796);
	nand 	XG7498 	(II19619,II19618,WX5795);
	nand 	XG7499 	(II19612,II19611,WX5794);
	nand 	XG7500 	(II19605,II19604,WX5793);
	nand 	XG7501 	(II19598,II19597,WX5792);
	nand 	XG7502 	(II19591,II19590,WX5791);
	nand 	XG7503 	(II19584,II19583,WX5790);
	nand 	XG7504 	(II19577,II19576,WX5789);
	nand 	XG7505 	(II19570,II19569,WX5788);
	nand 	XG7506 	(II19563,II19562,WX5787);
	nand 	XG7507 	(II19556,II19555,WX5786);
	nand 	XG7508 	(II19549,II19548,WX5785);
	nand 	XG7509 	(II19542,II19541,WX5784);
	nand 	XG7510 	(II15530,II15529,WX4522);
	nand 	XG7511 	(II15726,II15725,WX4521);
	nand 	XG7512 	(II15719,II15718,WX4520);
	nand 	XG7513 	(II15712,II15711,WX4519);
	nand 	XG7514 	(II15516,II15515,WX4518);
	nand 	XG7515 	(II15705,II15704,WX4517);
	nand 	XG7516 	(II15698,II15697,WX4516);
	nand 	XG7517 	(II15691,II15690,WX4515);
	nand 	XG7518 	(II15684,II15683,WX4514);
	nand 	XG7519 	(II15677,II15676,WX4513);
	nand 	XG7520 	(II15670,II15669,WX4512);
	nand 	XG7521 	(II15501,II15500,WX4511);
	nand 	XG7522 	(II15663,II15662,WX4510);
	nand 	XG7523 	(II15656,II15655,WX4509);
	nand 	XG7524 	(II15649,II15648,WX4508);
	nand 	XG7525 	(II15642,II15641,WX4507);
	nand 	XG7526 	(II15486,II15485,WX4506);
	nand 	XG7527 	(II15635,II15634,WX4505);
	nand 	XG7528 	(II15628,II15627,WX4504);
	nand 	XG7529 	(II15621,II15620,WX4503);
	nand 	XG7530 	(II15614,II15613,WX4502);
	nand 	XG7531 	(II15607,II15606,WX4501);
	nand 	XG7532 	(II15600,II15599,WX4500);
	nand 	XG7533 	(II15593,II15592,WX4499);
	nand 	XG7534 	(II15586,II15585,WX4498);
	nand 	XG7535 	(II15579,II15578,WX4497);
	nand 	XG7536 	(II15572,II15571,WX4496);
	nand 	XG7537 	(II15565,II15564,WX4495);
	nand 	XG7538 	(II15558,II15557,WX4494);
	nand 	XG7539 	(II15551,II15550,WX4493);
	nand 	XG7540 	(II15544,II15543,WX4492);
	nand 	XG7541 	(II15537,II15536,WX4491);
	nand 	XG7542 	(II11525,II11524,WX3229);
	nand 	XG7543 	(II11721,II11720,WX3228);
	nand 	XG7544 	(II11714,II11713,WX3227);
	nand 	XG7545 	(II11707,II11706,WX3226);
	nand 	XG7546 	(II11511,II11510,WX3225);
	nand 	XG7547 	(II11700,II11699,WX3224);
	nand 	XG7548 	(II11693,II11692,WX3223);
	nand 	XG7549 	(II11686,II11685,WX3222);
	nand 	XG7550 	(II11679,II11678,WX3221);
	nand 	XG7551 	(II11672,II11671,WX3220);
	nand 	XG7552 	(II11665,II11664,WX3219);
	nand 	XG7553 	(II11496,II11495,WX3218);
	nand 	XG7554 	(II11658,II11657,WX3217);
	nand 	XG7555 	(II11651,II11650,WX3216);
	nand 	XG7556 	(II11644,II11643,WX3215);
	nand 	XG7557 	(II11637,II11636,WX3214);
	nand 	XG7558 	(II11481,II11480,WX3213);
	nand 	XG7559 	(II11630,II11629,WX3212);
	nand 	XG7560 	(II11623,II11622,WX3211);
	nand 	XG7561 	(II11616,II11615,WX3210);
	nand 	XG7562 	(II11609,II11608,WX3209);
	nand 	XG7563 	(II11602,II11601,WX3208);
	nand 	XG7564 	(II11595,II11594,WX3207);
	nand 	XG7565 	(II11588,II11587,WX3206);
	nand 	XG7566 	(II11581,II11580,WX3205);
	nand 	XG7567 	(II11574,II11573,WX3204);
	nand 	XG7568 	(II11567,II11566,WX3203);
	nand 	XG7569 	(II11560,II11559,WX3202);
	nand 	XG7570 	(II11553,II11552,WX3201);
	nand 	XG7571 	(II11546,II11545,WX3200);
	nand 	XG7572 	(II11539,II11538,WX3199);
	nand 	XG7573 	(II11532,II11531,WX3198);
	nand 	XG7574 	(II7520,II7519,WX1936);
	nand 	XG7575 	(II7716,II7715,WX1935);
	nand 	XG7576 	(II7709,II7708,WX1934);
	nand 	XG7577 	(II7702,II7701,WX1933);
	nand 	XG7578 	(II7506,II7505,WX1932);
	nand 	XG7579 	(II7695,II7694,WX1931);
	nand 	XG7580 	(II7688,II7687,WX1930);
	nand 	XG7581 	(II7681,II7680,WX1929);
	nand 	XG7582 	(II7674,II7673,WX1928);
	nand 	XG7583 	(II7667,II7666,WX1927);
	nand 	XG7584 	(II7660,II7659,WX1926);
	nand 	XG7585 	(II7491,II7490,WX1925);
	nand 	XG7586 	(II7653,II7652,WX1924);
	nand 	XG7587 	(II7646,II7645,WX1923);
	nand 	XG7588 	(II7639,II7638,WX1922);
	nand 	XG7589 	(II7632,II7631,WX1921);
	nand 	XG7590 	(II7476,II7475,WX1920);
	nand 	XG7591 	(II7625,II7624,WX1919);
	nand 	XG7592 	(II7618,II7617,WX1918);
	nand 	XG7593 	(II7611,II7610,WX1917);
	nand 	XG7594 	(II7604,II7603,WX1916);
	nand 	XG7595 	(II7597,II7596,WX1915);
	nand 	XG7596 	(II7590,II7589,WX1914);
	nand 	XG7597 	(II7583,II7582,WX1913);
	nand 	XG7598 	(II7576,II7575,WX1912);
	nand 	XG7599 	(II7569,II7568,WX1911);
	nand 	XG7600 	(II7562,II7561,WX1910);
	nand 	XG7601 	(II7555,II7554,WX1909);
	nand 	XG7602 	(II7548,II7547,WX1908);
	nand 	XG7603 	(II7541,II7540,WX1907);
	nand 	XG7604 	(II7534,II7533,WX1906);
	nand 	XG7605 	(II7527,II7526,WX1905);
	nand 	XG7606 	(II3515,II3514,WX643);
	nand 	XG7607 	(II3711,II3710,WX642);
	nand 	XG7608 	(II3704,II3703,WX641);
	nand 	XG7609 	(II3697,II3696,WX640);
	nand 	XG7610 	(II3501,II3500,WX639);
	nand 	XG7611 	(II3690,II3689,WX638);
	nand 	XG7612 	(II3683,II3682,WX637);
	nand 	XG7613 	(II3676,II3675,WX636);
	nand 	XG7614 	(II3669,II3668,WX635);
	nand 	XG7615 	(II3662,II3661,WX634);
	nand 	XG7616 	(II3655,II3654,WX633);
	nand 	XG7617 	(II3486,II3485,WX632);
	nand 	XG7618 	(II3648,II3647,WX631);
	nand 	XG7619 	(II3641,II3640,WX630);
	nand 	XG7620 	(II3634,II3633,WX629);
	nand 	XG7621 	(II3627,II3626,WX628);
	nand 	XG7622 	(II3471,II3470,WX627);
	nand 	XG7623 	(II3620,II3619,WX626);
	nand 	XG7624 	(II3613,II3612,WX625);
	nand 	XG7625 	(II3606,II3605,WX624);
	nand 	XG7626 	(II3599,II3598,WX623);
	nand 	XG7627 	(II3592,II3591,WX622);
	nand 	XG7628 	(II3585,II3584,WX621);
	nand 	XG7629 	(II3578,II3577,WX620);
	nand 	XG7630 	(II3571,II3570,WX619);
	nand 	XG7631 	(II3564,II3563,WX618);
	nand 	XG7632 	(II3557,II3556,WX617);
	nand 	XG7633 	(II3550,II3549,WX616);
	nand 	XG7634 	(II3543,II3542,WX615);
	nand 	XG7635 	(II3536,II3535,WX614);
	nand 	XG7636 	(II3529,II3528,WX613);
	nand 	XG7637 	(II3522,II3521,WX612);
	nand 	XG7638 	(II3712,II3710,CRC_OUT_9_0);
	nand 	XG7639 	(II3705,II3703,CRC_OUT_9_1);
	nand 	XG7640 	(II3698,II3696,CRC_OUT_9_2);
	nand 	XG7641 	(II3691,II3689,CRC_OUT_9_4);
	nand 	XG7642 	(II3684,II3682,CRC_OUT_9_5);
	nand 	XG7643 	(II3677,II3675,CRC_OUT_9_6);
	nand 	XG7644 	(II3670,II3668,CRC_OUT_9_7);
	nand 	XG7645 	(II3663,II3661,CRC_OUT_9_8);
	nand 	XG7646 	(II3656,II3654,CRC_OUT_9_9);
	nand 	XG7647 	(II3649,II3647,CRC_OUT_9_11);
	nand 	XG7648 	(II3642,II3640,CRC_OUT_9_12);
	nand 	XG7649 	(II3635,II3633,CRC_OUT_9_13);
	nand 	XG7650 	(II3628,II3626,CRC_OUT_9_14);
	nand 	XG7651 	(II3621,II3619,CRC_OUT_9_16);
	nand 	XG7652 	(II3614,II3612,CRC_OUT_9_17);
	nand 	XG7653 	(II3607,II3605,CRC_OUT_9_18);
	nand 	XG7654 	(II3600,II3598,CRC_OUT_9_19);
	nand 	XG7655 	(II3593,II3591,CRC_OUT_9_20);
	nand 	XG7656 	(II3586,II3584,CRC_OUT_9_21);
	nand 	XG7657 	(II3579,II3577,CRC_OUT_9_22);
	nand 	XG7658 	(II3572,II3570,CRC_OUT_9_23);
	nand 	XG7659 	(II3565,II3563,CRC_OUT_9_24);
	nand 	XG7660 	(II3558,II3556,CRC_OUT_9_25);
	nand 	XG7661 	(II3551,II3549,CRC_OUT_9_26);
	nand 	XG7662 	(II3544,II3542,CRC_OUT_9_27);
	nand 	XG7663 	(II3537,II3535,CRC_OUT_9_28);
	nand 	XG7664 	(II3530,II3528,CRC_OUT_9_29);
	nand 	XG7665 	(II3523,II3521,CRC_OUT_9_30);
	nand 	XG7666 	(II3516,II3514,CRC_OUT_9_31);
	nand 	XG7667 	(II3502,II3500,CRC_OUT_9_31);
	nand 	XG7668 	(II3487,II3485,CRC_OUT_9_31);
	nand 	XG7669 	(II3472,II3470,CRC_OUT_9_31);
	nand 	XG7670 	(II7717,II7715,CRC_OUT_8_0);
	nand 	XG7671 	(II7710,II7708,CRC_OUT_8_1);
	nand 	XG7672 	(II7703,II7701,CRC_OUT_8_2);
	nand 	XG7673 	(II7696,II7694,CRC_OUT_8_4);
	nand 	XG7674 	(II7689,II7687,CRC_OUT_8_5);
	nand 	XG7675 	(II7682,II7680,CRC_OUT_8_6);
	nand 	XG7676 	(II7675,II7673,CRC_OUT_8_7);
	nand 	XG7677 	(II7668,II7666,CRC_OUT_8_8);
	nand 	XG7678 	(II7661,II7659,CRC_OUT_8_9);
	nand 	XG7679 	(II7654,II7652,CRC_OUT_8_11);
	nand 	XG7680 	(II7647,II7645,CRC_OUT_8_12);
	nand 	XG7681 	(II7640,II7638,CRC_OUT_8_13);
	nand 	XG7682 	(II7633,II7631,CRC_OUT_8_14);
	nand 	XG7683 	(II7626,II7624,CRC_OUT_8_16);
	nand 	XG7684 	(II7619,II7617,CRC_OUT_8_17);
	nand 	XG7685 	(II7612,II7610,CRC_OUT_8_18);
	nand 	XG7686 	(II7605,II7603,CRC_OUT_8_19);
	nand 	XG7687 	(II7598,II7596,CRC_OUT_8_20);
	nand 	XG7688 	(II7591,II7589,CRC_OUT_8_21);
	nand 	XG7689 	(II7584,II7582,CRC_OUT_8_22);
	nand 	XG7690 	(II7577,II7575,CRC_OUT_8_23);
	nand 	XG7691 	(II7570,II7568,CRC_OUT_8_24);
	nand 	XG7692 	(II7563,II7561,CRC_OUT_8_25);
	nand 	XG7693 	(II7556,II7554,CRC_OUT_8_26);
	nand 	XG7694 	(II7549,II7547,CRC_OUT_8_27);
	nand 	XG7695 	(II7542,II7540,CRC_OUT_8_28);
	nand 	XG7696 	(II7535,II7533,CRC_OUT_8_29);
	nand 	XG7697 	(II7528,II7526,CRC_OUT_8_30);
	nand 	XG7698 	(II7521,II7519,CRC_OUT_8_31);
	nand 	XG7699 	(II7507,II7505,CRC_OUT_8_31);
	nand 	XG7700 	(II7492,II7490,CRC_OUT_8_31);
	nand 	XG7701 	(II7477,II7475,CRC_OUT_8_31);
	nand 	XG7702 	(II11722,II11720,CRC_OUT_7_0);
	nand 	XG7703 	(II11715,II11713,CRC_OUT_7_1);
	nand 	XG7704 	(II11708,II11706,CRC_OUT_7_2);
	nand 	XG7705 	(II11701,II11699,CRC_OUT_7_4);
	nand 	XG7706 	(II11694,II11692,CRC_OUT_7_5);
	nand 	XG7707 	(II11687,II11685,CRC_OUT_7_6);
	nand 	XG7708 	(II11680,II11678,CRC_OUT_7_7);
	nand 	XG7709 	(II11673,II11671,CRC_OUT_7_8);
	nand 	XG7710 	(II11666,II11664,CRC_OUT_7_9);
	nand 	XG7711 	(II11659,II11657,CRC_OUT_7_11);
	nand 	XG7712 	(II11652,II11650,CRC_OUT_7_12);
	nand 	XG7713 	(II11645,II11643,CRC_OUT_7_13);
	nand 	XG7714 	(II11638,II11636,CRC_OUT_7_14);
	nand 	XG7715 	(II11631,II11629,CRC_OUT_7_16);
	nand 	XG7716 	(II11624,II11622,CRC_OUT_7_17);
	nand 	XG7717 	(II11617,II11615,CRC_OUT_7_18);
	nand 	XG7718 	(II11610,II11608,CRC_OUT_7_19);
	nand 	XG7719 	(II11603,II11601,CRC_OUT_7_20);
	nand 	XG7720 	(II11596,II11594,CRC_OUT_7_21);
	nand 	XG7721 	(II11589,II11587,CRC_OUT_7_22);
	nand 	XG7722 	(II11582,II11580,CRC_OUT_7_23);
	nand 	XG7723 	(II11575,II11573,CRC_OUT_7_24);
	nand 	XG7724 	(II11568,II11566,CRC_OUT_7_25);
	nand 	XG7725 	(II11561,II11559,CRC_OUT_7_26);
	nand 	XG7726 	(II11554,II11552,CRC_OUT_7_27);
	nand 	XG7727 	(II11547,II11545,CRC_OUT_7_28);
	nand 	XG7728 	(II11540,II11538,CRC_OUT_7_29);
	nand 	XG7729 	(II11533,II11531,CRC_OUT_7_30);
	nand 	XG7730 	(II11526,II11524,CRC_OUT_7_31);
	nand 	XG7731 	(II11512,II11510,CRC_OUT_7_31);
	nand 	XG7732 	(II11497,II11495,CRC_OUT_7_31);
	nand 	XG7733 	(II11482,II11480,CRC_OUT_7_31);
	nand 	XG7734 	(II15727,II15725,CRC_OUT_6_0);
	nand 	XG7735 	(II15720,II15718,CRC_OUT_6_1);
	nand 	XG7736 	(II15713,II15711,CRC_OUT_6_2);
	nand 	XG7737 	(II15706,II15704,CRC_OUT_6_4);
	nand 	XG7738 	(II15699,II15697,CRC_OUT_6_5);
	nand 	XG7739 	(II15692,II15690,CRC_OUT_6_6);
	nand 	XG7740 	(II15685,II15683,CRC_OUT_6_7);
	nand 	XG7741 	(II15678,II15676,CRC_OUT_6_8);
	nand 	XG7742 	(II15671,II15669,CRC_OUT_6_9);
	nand 	XG7743 	(II15664,II15662,CRC_OUT_6_11);
	nand 	XG7744 	(II15657,II15655,CRC_OUT_6_12);
	nand 	XG7745 	(II15650,II15648,CRC_OUT_6_13);
	nand 	XG7746 	(II15643,II15641,CRC_OUT_6_14);
	nand 	XG7747 	(II15636,II15634,CRC_OUT_6_16);
	nand 	XG7748 	(II15629,II15627,CRC_OUT_6_17);
	nand 	XG7749 	(II15622,II15620,CRC_OUT_6_18);
	nand 	XG7750 	(II15615,II15613,CRC_OUT_6_19);
	nand 	XG7751 	(II15608,II15606,CRC_OUT_6_20);
	nand 	XG7752 	(II15601,II15599,CRC_OUT_6_21);
	nand 	XG7753 	(II15594,II15592,CRC_OUT_6_22);
	nand 	XG7754 	(II15587,II15585,CRC_OUT_6_23);
	nand 	XG7755 	(II15580,II15578,CRC_OUT_6_24);
	nand 	XG7756 	(II15573,II15571,CRC_OUT_6_25);
	nand 	XG7757 	(II15566,II15564,CRC_OUT_6_26);
	nand 	XG7758 	(II15559,II15557,CRC_OUT_6_27);
	nand 	XG7759 	(II15552,II15550,CRC_OUT_6_28);
	nand 	XG7760 	(II15545,II15543,CRC_OUT_6_29);
	nand 	XG7761 	(II15538,II15536,CRC_OUT_6_30);
	nand 	XG7762 	(II15531,II15529,CRC_OUT_6_31);
	nand 	XG7763 	(II15517,II15515,CRC_OUT_6_31);
	nand 	XG7764 	(II15502,II15500,CRC_OUT_6_31);
	nand 	XG7765 	(II15487,II15485,CRC_OUT_6_31);
	nand 	XG7766 	(II19732,II19730,CRC_OUT_5_0);
	nand 	XG7767 	(II19725,II19723,CRC_OUT_5_1);
	nand 	XG7768 	(II19718,II19716,CRC_OUT_5_2);
	nand 	XG7769 	(II19711,II19709,CRC_OUT_5_4);
	nand 	XG7770 	(II19704,II19702,CRC_OUT_5_5);
	nand 	XG7771 	(II19697,II19695,CRC_OUT_5_6);
	nand 	XG7772 	(II19690,II19688,CRC_OUT_5_7);
	nand 	XG7773 	(II19683,II19681,CRC_OUT_5_8);
	nand 	XG7774 	(II19676,II19674,CRC_OUT_5_9);
	nand 	XG7775 	(II19669,II19667,CRC_OUT_5_11);
	nand 	XG7776 	(II19662,II19660,CRC_OUT_5_12);
	nand 	XG7777 	(II19655,II19653,CRC_OUT_5_13);
	nand 	XG7778 	(II19648,II19646,CRC_OUT_5_14);
	nand 	XG7779 	(II19641,II19639,CRC_OUT_5_16);
	nand 	XG7780 	(II19634,II19632,CRC_OUT_5_17);
	nand 	XG7781 	(II19627,II19625,CRC_OUT_5_18);
	nand 	XG7782 	(II19620,II19618,CRC_OUT_5_19);
	nand 	XG7783 	(II19613,II19611,CRC_OUT_5_20);
	nand 	XG7784 	(II19606,II19604,CRC_OUT_5_21);
	nand 	XG7785 	(II19599,II19597,CRC_OUT_5_22);
	nand 	XG7786 	(II19592,II19590,CRC_OUT_5_23);
	nand 	XG7787 	(II19585,II19583,CRC_OUT_5_24);
	nand 	XG7788 	(II19578,II19576,CRC_OUT_5_25);
	nand 	XG7789 	(II19571,II19569,CRC_OUT_5_26);
	nand 	XG7790 	(II19564,II19562,CRC_OUT_5_27);
	nand 	XG7791 	(II19557,II19555,CRC_OUT_5_28);
	nand 	XG7792 	(II19550,II19548,CRC_OUT_5_29);
	nand 	XG7793 	(II19543,II19541,CRC_OUT_5_30);
	nand 	XG7794 	(II19536,II19534,CRC_OUT_5_31);
	nand 	XG7795 	(II19522,II19520,CRC_OUT_5_31);
	nand 	XG7796 	(II19507,II19505,CRC_OUT_5_31);
	nand 	XG7797 	(II19492,II19490,CRC_OUT_5_31);
	nand 	XG7798 	(II23737,II23735,CRC_OUT_4_0);
	nand 	XG7799 	(II23730,II23728,CRC_OUT_4_1);
	nand 	XG7800 	(II23723,II23721,CRC_OUT_4_2);
	nand 	XG7801 	(II23716,II23714,CRC_OUT_4_4);
	nand 	XG7802 	(II23709,II23707,CRC_OUT_4_5);
	nand 	XG7803 	(II23702,II23700,CRC_OUT_4_6);
	nand 	XG7804 	(II23695,II23693,CRC_OUT_4_7);
	nand 	XG7805 	(II23688,II23686,CRC_OUT_4_8);
	nand 	XG7806 	(II23681,II23679,CRC_OUT_4_9);
	nand 	XG7807 	(II23674,II23672,CRC_OUT_4_11);
	nand 	XG7808 	(II23667,II23665,CRC_OUT_4_12);
	nand 	XG7809 	(II23660,II23658,CRC_OUT_4_13);
	nand 	XG7810 	(II23653,II23651,CRC_OUT_4_14);
	nand 	XG7811 	(II23646,II23644,CRC_OUT_4_16);
	nand 	XG7812 	(II23639,II23637,CRC_OUT_4_17);
	nand 	XG7813 	(II23632,II23630,CRC_OUT_4_18);
	nand 	XG7814 	(II23625,II23623,CRC_OUT_4_19);
	nand 	XG7815 	(II23618,II23616,CRC_OUT_4_20);
	nand 	XG7816 	(II23611,II23609,CRC_OUT_4_21);
	nand 	XG7817 	(II23604,II23602,CRC_OUT_4_22);
	nand 	XG7818 	(II23597,II23595,CRC_OUT_4_23);
	nand 	XG7819 	(II23590,II23588,CRC_OUT_4_24);
	nand 	XG7820 	(II23583,II23581,CRC_OUT_4_25);
	nand 	XG7821 	(II23576,II23574,CRC_OUT_4_26);
	nand 	XG7822 	(II23569,II23567,CRC_OUT_4_27);
	nand 	XG7823 	(II23562,II23560,CRC_OUT_4_28);
	nand 	XG7824 	(II23555,II23553,CRC_OUT_4_29);
	nand 	XG7825 	(II23548,II23546,CRC_OUT_4_30);
	nand 	XG7826 	(II23541,II23539,CRC_OUT_4_31);
	nand 	XG7827 	(II23527,II23525,CRC_OUT_4_31);
	nand 	XG7828 	(II23512,II23510,CRC_OUT_4_31);
	nand 	XG7829 	(II23497,II23495,CRC_OUT_4_31);
	nand 	XG7830 	(II27742,II27740,CRC_OUT_3_0);
	nand 	XG7831 	(II27735,II27733,CRC_OUT_3_1);
	nand 	XG7832 	(II27728,II27726,CRC_OUT_3_2);
	nand 	XG7833 	(II27721,II27719,CRC_OUT_3_4);
	nand 	XG7834 	(II27714,II27712,CRC_OUT_3_5);
	nand 	XG7835 	(II27707,II27705,CRC_OUT_3_6);
	nand 	XG7836 	(II27700,II27698,CRC_OUT_3_7);
	nand 	XG7837 	(II27693,II27691,CRC_OUT_3_8);
	nand 	XG7838 	(II27686,II27684,CRC_OUT_3_9);
	nand 	XG7839 	(II27679,II27677,CRC_OUT_3_11);
	nand 	XG7840 	(II27672,II27670,CRC_OUT_3_12);
	nand 	XG7841 	(II27665,II27663,CRC_OUT_3_13);
	nand 	XG7842 	(II27658,II27656,CRC_OUT_3_14);
	nand 	XG7843 	(II27651,II27649,CRC_OUT_3_16);
	nand 	XG7844 	(II27644,II27642,CRC_OUT_3_17);
	nand 	XG7845 	(II27637,II27635,CRC_OUT_3_18);
	nand 	XG7846 	(II27630,II27628,CRC_OUT_3_19);
	nand 	XG7847 	(II27623,II27621,CRC_OUT_3_20);
	nand 	XG7848 	(II27616,II27614,CRC_OUT_3_21);
	nand 	XG7849 	(II27609,II27607,CRC_OUT_3_22);
	nand 	XG7850 	(II27602,II27600,CRC_OUT_3_23);
	nand 	XG7851 	(II27595,II27593,CRC_OUT_3_24);
	nand 	XG7852 	(II27588,II27586,CRC_OUT_3_25);
	nand 	XG7853 	(II27581,II27579,CRC_OUT_3_26);
	nand 	XG7854 	(II27574,II27572,CRC_OUT_3_27);
	nand 	XG7855 	(II27567,II27565,CRC_OUT_3_28);
	nand 	XG7856 	(II27560,II27558,CRC_OUT_3_29);
	nand 	XG7857 	(II27553,II27551,CRC_OUT_3_30);
	nand 	XG7858 	(II27546,II27544,CRC_OUT_3_31);
	nand 	XG7859 	(II27532,II27530,CRC_OUT_3_31);
	nand 	XG7860 	(II27517,II27515,CRC_OUT_3_31);
	nand 	XG7861 	(II27502,II27500,CRC_OUT_3_31);
	nand 	XG7862 	(II31747,II31745,CRC_OUT_2_0);
	nand 	XG7863 	(II31740,II31738,CRC_OUT_2_1);
	nand 	XG7864 	(II31733,II31731,CRC_OUT_2_2);
	nand 	XG7865 	(II31726,II31724,CRC_OUT_2_4);
	nand 	XG7866 	(II31719,II31717,CRC_OUT_2_5);
	nand 	XG7867 	(II31712,II31710,CRC_OUT_2_6);
	nand 	XG7868 	(II31705,II31703,CRC_OUT_2_7);
	nand 	XG7869 	(II31698,II31696,CRC_OUT_2_8);
	nand 	XG7870 	(II31691,II31689,CRC_OUT_2_9);
	nand 	XG7871 	(II31684,II31682,CRC_OUT_2_11);
	nand 	XG7872 	(II31677,II31675,CRC_OUT_2_12);
	nand 	XG7873 	(II31670,II31668,CRC_OUT_2_13);
	nand 	XG7874 	(II31663,II31661,CRC_OUT_2_14);
	nand 	XG7875 	(II31656,II31654,CRC_OUT_2_16);
	nand 	XG7876 	(II31649,II31647,CRC_OUT_2_17);
	nand 	XG7877 	(II31642,II31640,CRC_OUT_2_18);
	nand 	XG7878 	(II31635,II31633,CRC_OUT_2_19);
	nand 	XG7879 	(II31628,II31626,CRC_OUT_2_20);
	nand 	XG7880 	(II31621,II31619,CRC_OUT_2_21);
	nand 	XG7881 	(II31614,II31612,CRC_OUT_2_22);
	nand 	XG7882 	(II31607,II31605,CRC_OUT_2_23);
	nand 	XG7883 	(II31600,II31598,CRC_OUT_2_24);
	nand 	XG7884 	(II31593,II31591,CRC_OUT_2_25);
	nand 	XG7885 	(II31586,II31584,CRC_OUT_2_26);
	nand 	XG7886 	(II31579,II31577,CRC_OUT_2_27);
	nand 	XG7887 	(II31572,II31570,CRC_OUT_2_28);
	nand 	XG7888 	(II31565,II31563,CRC_OUT_2_29);
	nand 	XG7889 	(II31558,II31556,CRC_OUT_2_30);
	nand 	XG7890 	(II31551,II31549,CRC_OUT_2_31);
	nand 	XG7891 	(II31537,II31535,CRC_OUT_2_31);
	nand 	XG7892 	(II31522,II31520,CRC_OUT_2_31);
	nand 	XG7893 	(II31507,II31505,CRC_OUT_2_31);
	nand 	XG7894 	(II35752,II35750,CRC_OUT_1_0);
	nand 	XG7895 	(II35745,II35743,CRC_OUT_1_1);
	nand 	XG7896 	(II35738,II35736,CRC_OUT_1_2);
	nand 	XG7897 	(II35731,II35729,CRC_OUT_1_4);
	nand 	XG7898 	(II35724,II35722,CRC_OUT_1_5);
	nand 	XG7899 	(II35717,II35715,CRC_OUT_1_6);
	nand 	XG7900 	(II35710,II35708,CRC_OUT_1_7);
	nand 	XG7901 	(II35703,II35701,CRC_OUT_1_8);
	nand 	XG7902 	(II35696,II35694,CRC_OUT_1_9);
	nand 	XG7903 	(II35689,II35687,CRC_OUT_1_11);
	nand 	XG7904 	(II35682,II35680,CRC_OUT_1_12);
	nand 	XG7905 	(II35675,II35673,CRC_OUT_1_13);
	nand 	XG7906 	(II35668,II35666,CRC_OUT_1_14);
	nand 	XG7907 	(II35661,II35659,CRC_OUT_1_16);
	nand 	XG7908 	(II35654,II35652,CRC_OUT_1_17);
	nand 	XG7909 	(II35647,II35645,CRC_OUT_1_18);
	nand 	XG7910 	(II35640,II35638,CRC_OUT_1_19);
	nand 	XG7911 	(II35633,II35631,CRC_OUT_1_20);
	nand 	XG7912 	(II35626,II35624,CRC_OUT_1_21);
	nand 	XG7913 	(II35619,II35617,CRC_OUT_1_22);
	nand 	XG7914 	(II35612,II35610,CRC_OUT_1_23);
	nand 	XG7915 	(II35605,II35603,CRC_OUT_1_24);
	nand 	XG7916 	(II35598,II35596,CRC_OUT_1_25);
	nand 	XG7917 	(II35591,II35589,CRC_OUT_1_26);
	nand 	XG7918 	(II35584,II35582,CRC_OUT_1_27);
	nand 	XG7919 	(II35577,II35575,CRC_OUT_1_28);
	nand 	XG7920 	(II35570,II35568,CRC_OUT_1_29);
	nand 	XG7921 	(II35563,II35561,CRC_OUT_1_30);
	nand 	XG7922 	(II35556,II35554,CRC_OUT_1_31);
	nand 	XG7923 	(II35542,II35540,CRC_OUT_1_31);
	nand 	XG7924 	(II35527,II35525,CRC_OUT_1_31);
	nand 	XG7925 	(II35512,II35510,CRC_OUT_1_31);
	nand 	XG7926 	(II34988,II34991,II34990);
	nand 	XG7927 	(II34957,II34960,II34959);
	nand 	XG7928 	(II34926,II34929,II34928);
	nand 	XG7929 	(II34895,II34898,II34897);
	nand 	XG7930 	(II34864,II34867,II34866);
	nand 	XG7931 	(II34833,II34836,II34835);
	nand 	XG7932 	(II34802,II34805,II34804);
	nand 	XG7933 	(II34771,II34774,II34773);
	nand 	XG7934 	(II34740,II34743,II34742);
	nand 	XG7935 	(II34709,II34712,II34711);
	nand 	XG7936 	(II34678,II34681,II34680);
	nand 	XG7937 	(II34647,II34650,II34649);
	nand 	XG7938 	(II34616,II34619,II34618);
	nand 	XG7939 	(II34585,II34588,II34587);
	nand 	XG7940 	(II34554,II34557,II34556);
	nand 	XG7941 	(II34523,II34526,II34525);
	nand 	XG7942 	(II34492,II34495,II34494);
	nand 	XG7943 	(II34461,II34464,II34463);
	nand 	XG7944 	(II34430,II34433,II34432);
	nand 	XG7945 	(II34399,II34402,II34401);
	nand 	XG7946 	(II34368,II34371,II34370);
	nand 	XG7947 	(II34337,II34340,II34339);
	nand 	XG7948 	(II34306,II34309,II34308);
	nand 	XG7949 	(II34275,II34278,II34277);
	nand 	XG7950 	(II34244,II34247,II34246);
	nand 	XG7951 	(II34213,II34216,II34215);
	nand 	XG7952 	(II34182,II34185,II34184);
	nand 	XG7953 	(II34151,II34154,II34153);
	nand 	XG7954 	(II34120,II34123,II34122);
	nand 	XG7955 	(II34089,II34092,II34091);
	nand 	XG7956 	(II34058,II34061,II34060);
	nand 	XG7957 	(II34027,II34030,II34029);
	nand 	XG7958 	(II30983,II30986,II30985);
	nand 	XG7959 	(II30952,II30955,II30954);
	nand 	XG7960 	(II30921,II30924,II30923);
	nand 	XG7961 	(II30890,II30893,II30892);
	nand 	XG7962 	(II30859,II30862,II30861);
	nand 	XG7963 	(II30828,II30831,II30830);
	nand 	XG7964 	(II30797,II30800,II30799);
	nand 	XG7965 	(II30766,II30769,II30768);
	nand 	XG7966 	(II30735,II30738,II30737);
	nand 	XG7967 	(II30704,II30707,II30706);
	nand 	XG7968 	(II30673,II30676,II30675);
	nand 	XG7969 	(II30642,II30645,II30644);
	nand 	XG7970 	(II30611,II30614,II30613);
	nand 	XG7971 	(II30580,II30583,II30582);
	nand 	XG7972 	(II30549,II30552,II30551);
	nand 	XG7973 	(II30518,II30521,II30520);
	nand 	XG7974 	(II30487,II30490,II30489);
	nand 	XG7975 	(II30456,II30459,II30458);
	nand 	XG7976 	(II30425,II30428,II30427);
	nand 	XG7977 	(II30394,II30397,II30396);
	nand 	XG7978 	(II30363,II30366,II30365);
	nand 	XG7979 	(II30332,II30335,II30334);
	nand 	XG7980 	(II30301,II30304,II30303);
	nand 	XG7981 	(II30270,II30273,II30272);
	nand 	XG7982 	(II30239,II30242,II30241);
	nand 	XG7983 	(II30208,II30211,II30210);
	nand 	XG7984 	(II30177,II30180,II30179);
	nand 	XG7985 	(II30146,II30149,II30148);
	nand 	XG7986 	(II30115,II30118,II30117);
	nand 	XG7987 	(II30084,II30087,II30086);
	nand 	XG7988 	(II30053,II30056,II30055);
	nand 	XG7989 	(II30022,II30025,II30024);
	nand 	XG7990 	(II26978,II26981,II26980);
	nand 	XG7991 	(II26947,II26950,II26949);
	nand 	XG7992 	(II26916,II26919,II26918);
	nand 	XG7993 	(II26885,II26888,II26887);
	nand 	XG7994 	(II26854,II26857,II26856);
	nand 	XG7995 	(II26823,II26826,II26825);
	nand 	XG7996 	(II26792,II26795,II26794);
	nand 	XG7997 	(II26761,II26764,II26763);
	nand 	XG7998 	(II26730,II26733,II26732);
	nand 	XG7999 	(II26699,II26702,II26701);
	nand 	XG8000 	(II26668,II26671,II26670);
	nand 	XG8001 	(II26637,II26640,II26639);
	nand 	XG8002 	(II26606,II26609,II26608);
	nand 	XG8003 	(II26575,II26578,II26577);
	nand 	XG8004 	(II26544,II26547,II26546);
	nand 	XG8005 	(II26513,II26516,II26515);
	nand 	XG8006 	(II26482,II26485,II26484);
	nand 	XG8007 	(II26451,II26454,II26453);
	nand 	XG8008 	(II26420,II26423,II26422);
	nand 	XG8009 	(II26389,II26392,II26391);
	nand 	XG8010 	(II26358,II26361,II26360);
	nand 	XG8011 	(II26327,II26330,II26329);
	nand 	XG8012 	(II26296,II26299,II26298);
	nand 	XG8013 	(II26265,II26268,II26267);
	nand 	XG8014 	(II26234,II26237,II26236);
	nand 	XG8015 	(II26203,II26206,II26205);
	nand 	XG8016 	(II26172,II26175,II26174);
	nand 	XG8017 	(II26141,II26144,II26143);
	nand 	XG8018 	(II26110,II26113,II26112);
	nand 	XG8019 	(II26079,II26082,II26081);
	nand 	XG8020 	(II26048,II26051,II26050);
	nand 	XG8021 	(II26017,II26020,II26019);
	nand 	XG8022 	(II22973,II22976,II22975);
	nand 	XG8023 	(II22942,II22945,II22944);
	nand 	XG8024 	(II22911,II22914,II22913);
	nand 	XG8025 	(II22880,II22883,II22882);
	nand 	XG8026 	(II22849,II22852,II22851);
	nand 	XG8027 	(II22818,II22821,II22820);
	nand 	XG8028 	(II22787,II22790,II22789);
	nand 	XG8029 	(II22756,II22759,II22758);
	nand 	XG8030 	(II22725,II22728,II22727);
	nand 	XG8031 	(II22694,II22697,II22696);
	nand 	XG8032 	(II22663,II22666,II22665);
	nand 	XG8033 	(II22632,II22635,II22634);
	nand 	XG8034 	(II22601,II22604,II22603);
	nand 	XG8035 	(II22570,II22573,II22572);
	nand 	XG8036 	(II22539,II22542,II22541);
	nand 	XG8037 	(II22508,II22511,II22510);
	nand 	XG8038 	(II22477,II22480,II22479);
	nand 	XG8039 	(II22446,II22449,II22448);
	nand 	XG8040 	(II22415,II22418,II22417);
	nand 	XG8041 	(II22384,II22387,II22386);
	nand 	XG8042 	(II22353,II22356,II22355);
	nand 	XG8043 	(II22322,II22325,II22324);
	nand 	XG8044 	(II22291,II22294,II22293);
	nand 	XG8045 	(II22260,II22263,II22262);
	nand 	XG8046 	(II22229,II22232,II22231);
	nand 	XG8047 	(II22198,II22201,II22200);
	nand 	XG8048 	(II22167,II22170,II22169);
	nand 	XG8049 	(II22136,II22139,II22138);
	nand 	XG8050 	(II22105,II22108,II22107);
	nand 	XG8051 	(II22074,II22077,II22076);
	nand 	XG8052 	(II22043,II22046,II22045);
	nand 	XG8053 	(II22012,II22015,II22014);
	nand 	XG8054 	(II18968,II18971,II18970);
	nand 	XG8055 	(II18937,II18940,II18939);
	nand 	XG8056 	(II18906,II18909,II18908);
	nand 	XG8057 	(II18875,II18878,II18877);
	nand 	XG8058 	(II18844,II18847,II18846);
	nand 	XG8059 	(II18813,II18816,II18815);
	nand 	XG8060 	(II18782,II18785,II18784);
	nand 	XG8061 	(II18751,II18754,II18753);
	nand 	XG8062 	(II18720,II18723,II18722);
	nand 	XG8063 	(II18689,II18692,II18691);
	nand 	XG8064 	(II18658,II18661,II18660);
	nand 	XG8065 	(II18627,II18630,II18629);
	nand 	XG8066 	(II18596,II18599,II18598);
	nand 	XG8067 	(II18565,II18568,II18567);
	nand 	XG8068 	(II18534,II18537,II18536);
	nand 	XG8069 	(II18503,II18506,II18505);
	nand 	XG8070 	(II18472,II18475,II18474);
	nand 	XG8071 	(II18441,II18444,II18443);
	nand 	XG8072 	(II18410,II18413,II18412);
	nand 	XG8073 	(II18379,II18382,II18381);
	nand 	XG8074 	(II18348,II18351,II18350);
	nand 	XG8075 	(II18317,II18320,II18319);
	nand 	XG8076 	(II18286,II18289,II18288);
	nand 	XG8077 	(II18255,II18258,II18257);
	nand 	XG8078 	(II18224,II18227,II18226);
	nand 	XG8079 	(II18193,II18196,II18195);
	nand 	XG8080 	(II18162,II18165,II18164);
	nand 	XG8081 	(II18131,II18134,II18133);
	nand 	XG8082 	(II18100,II18103,II18102);
	nand 	XG8083 	(II18069,II18072,II18071);
	nand 	XG8084 	(II18038,II18041,II18040);
	nand 	XG8085 	(II18007,II18010,II18009);
	nand 	XG8086 	(II14963,II14966,II14965);
	nand 	XG8087 	(II14932,II14935,II14934);
	nand 	XG8088 	(II14901,II14904,II14903);
	nand 	XG8089 	(II14870,II14873,II14872);
	nand 	XG8090 	(II14839,II14842,II14841);
	nand 	XG8091 	(II14808,II14811,II14810);
	nand 	XG8092 	(II14777,II14780,II14779);
	nand 	XG8093 	(II14746,II14749,II14748);
	nand 	XG8094 	(II14715,II14718,II14717);
	nand 	XG8095 	(II14684,II14687,II14686);
	nand 	XG8096 	(II14653,II14656,II14655);
	nand 	XG8097 	(II14622,II14625,II14624);
	nand 	XG8098 	(II14591,II14594,II14593);
	nand 	XG8099 	(II14560,II14563,II14562);
	nand 	XG8100 	(II14529,II14532,II14531);
	nand 	XG8101 	(II14498,II14501,II14500);
	nand 	XG8102 	(II14467,II14470,II14469);
	nand 	XG8103 	(II14436,II14439,II14438);
	nand 	XG8104 	(II14405,II14408,II14407);
	nand 	XG8105 	(II14374,II14377,II14376);
	nand 	XG8106 	(II14343,II14346,II14345);
	nand 	XG8107 	(II14312,II14315,II14314);
	nand 	XG8108 	(II14281,II14284,II14283);
	nand 	XG8109 	(II14250,II14253,II14252);
	nand 	XG8110 	(II14219,II14222,II14221);
	nand 	XG8111 	(II14188,II14191,II14190);
	nand 	XG8112 	(II14157,II14160,II14159);
	nand 	XG8113 	(II14126,II14129,II14128);
	nand 	XG8114 	(II14095,II14098,II14097);
	nand 	XG8115 	(II14064,II14067,II14066);
	nand 	XG8116 	(II14033,II14036,II14035);
	nand 	XG8117 	(II14002,II14005,II14004);
	nand 	XG8118 	(II10958,II10961,II10960);
	nand 	XG8119 	(II10927,II10930,II10929);
	nand 	XG8120 	(II10896,II10899,II10898);
	nand 	XG8121 	(II10865,II10868,II10867);
	nand 	XG8122 	(II10834,II10837,II10836);
	nand 	XG8123 	(II10803,II10806,II10805);
	nand 	XG8124 	(II10772,II10775,II10774);
	nand 	XG8125 	(II10741,II10744,II10743);
	nand 	XG8126 	(II10710,II10713,II10712);
	nand 	XG8127 	(II10679,II10682,II10681);
	nand 	XG8128 	(II10648,II10651,II10650);
	nand 	XG8129 	(II10617,II10620,II10619);
	nand 	XG8130 	(II10586,II10589,II10588);
	nand 	XG8131 	(II10555,II10558,II10557);
	nand 	XG8132 	(II10524,II10527,II10526);
	nand 	XG8133 	(II10493,II10496,II10495);
	nand 	XG8134 	(II10462,II10465,II10464);
	nand 	XG8135 	(II10431,II10434,II10433);
	nand 	XG8136 	(II10400,II10403,II10402);
	nand 	XG8137 	(II10369,II10372,II10371);
	nand 	XG8138 	(II10338,II10341,II10340);
	nand 	XG8139 	(II10307,II10310,II10309);
	nand 	XG8140 	(II10276,II10279,II10278);
	nand 	XG8141 	(II10245,II10248,II10247);
	nand 	XG8142 	(II10214,II10217,II10216);
	nand 	XG8143 	(II10183,II10186,II10185);
	nand 	XG8144 	(II10152,II10155,II10154);
	nand 	XG8145 	(II10121,II10124,II10123);
	nand 	XG8146 	(II10090,II10093,II10092);
	nand 	XG8147 	(II10059,II10062,II10061);
	nand 	XG8148 	(II10028,II10031,II10030);
	nand 	XG8149 	(II9997,II10000,II9999);
	nand 	XG8150 	(II6953,II6956,II6955);
	nand 	XG8151 	(II6922,II6925,II6924);
	nand 	XG8152 	(II6891,II6894,II6893);
	nand 	XG8153 	(II6860,II6863,II6862);
	nand 	XG8154 	(II6829,II6832,II6831);
	nand 	XG8155 	(II6798,II6801,II6800);
	nand 	XG8156 	(II6767,II6770,II6769);
	nand 	XG8157 	(II6736,II6739,II6738);
	nand 	XG8158 	(II6705,II6708,II6707);
	nand 	XG8159 	(II6674,II6677,II6676);
	nand 	XG8160 	(II6643,II6646,II6645);
	nand 	XG8161 	(II6612,II6615,II6614);
	nand 	XG8162 	(II6581,II6584,II6583);
	nand 	XG8163 	(II6550,II6553,II6552);
	nand 	XG8164 	(II6519,II6522,II6521);
	nand 	XG8165 	(II6488,II6491,II6490);
	nand 	XG8166 	(II6457,II6460,II6459);
	nand 	XG8167 	(II6426,II6429,II6428);
	nand 	XG8168 	(II6395,II6398,II6397);
	nand 	XG8169 	(II6364,II6367,II6366);
	nand 	XG8170 	(II6333,II6336,II6335);
	nand 	XG8171 	(II6302,II6305,II6304);
	nand 	XG8172 	(II6271,II6274,II6273);
	nand 	XG8173 	(II6240,II6243,II6242);
	nand 	XG8174 	(II6209,II6212,II6211);
	nand 	XG8175 	(II6178,II6181,II6180);
	nand 	XG8176 	(II6147,II6150,II6149);
	nand 	XG8177 	(II6116,II6119,II6118);
	nand 	XG8178 	(II6085,II6088,II6087);
	nand 	XG8179 	(II6054,II6057,II6056);
	nand 	XG8180 	(II6023,II6026,II6025);
	nand 	XG8181 	(II5992,II5995,II5994);
	nand 	XG8182 	(II2948,II2951,II2950);
	nand 	XG8183 	(II2917,II2920,II2919);
	nand 	XG8184 	(II2886,II2889,II2888);
	nand 	XG8185 	(II2855,II2858,II2857);
	nand 	XG8186 	(II2824,II2827,II2826);
	nand 	XG8187 	(II2793,II2796,II2795);
	nand 	XG8188 	(II2762,II2765,II2764);
	nand 	XG8189 	(II2731,II2734,II2733);
	nand 	XG8190 	(II2700,II2703,II2702);
	nand 	XG8191 	(II2669,II2672,II2671);
	nand 	XG8192 	(II2638,II2641,II2640);
	nand 	XG8193 	(II2607,II2610,II2609);
	nand 	XG8194 	(II2576,II2579,II2578);
	nand 	XG8195 	(II2545,II2548,II2547);
	nand 	XG8196 	(II2514,II2517,II2516);
	nand 	XG8197 	(II2483,II2486,II2485);
	nand 	XG8198 	(II2452,II2455,II2454);
	nand 	XG8199 	(II2421,II2424,II2423);
	nand 	XG8200 	(II2390,II2393,II2392);
	nand 	XG8201 	(II2359,II2362,II2361);
	nand 	XG8202 	(II2328,II2331,II2330);
	nand 	XG8203 	(II2297,II2300,II2299);
	nand 	XG8204 	(II2266,II2269,II2268);
	nand 	XG8205 	(II2235,II2238,II2237);
	nand 	XG8206 	(II2204,II2207,II2206);
	nand 	XG8207 	(II2173,II2176,II2175);
	nand 	XG8208 	(II2142,II2145,II2144);
	nand 	XG8209 	(II2111,II2114,II2113);
	nand 	XG8210 	(II2080,II2083,II2082);
	nand 	XG8211 	(II2049,II2052,II2051);
	nand 	XG8212 	(II2018,II2021,II2020);
	nand 	XG8213 	(II1987,II1990,II1989);
	or 	XG8214 	(WX10386,WX10383,WX10384);
	or 	XG8215 	(WX10400,WX10397,WX10398);
	or 	XG8216 	(WX10414,WX10411,WX10412);
	or 	XG8217 	(WX10428,WX10425,WX10426);
	or 	XG8218 	(WX10442,WX10439,WX10440);
	or 	XG8219 	(WX10456,WX10453,WX10454);
	or 	XG8220 	(WX10470,WX10467,WX10468);
	or 	XG8221 	(WX10484,WX10481,WX10482);
	or 	XG8222 	(WX10498,WX10495,WX10496);
	or 	XG8223 	(WX10512,WX10509,WX10510);
	or 	XG8224 	(WX10526,WX10523,WX10524);
	or 	XG8225 	(WX10540,WX10537,WX10538);
	or 	XG8226 	(WX10554,WX10551,WX10552);
	or 	XG8227 	(WX10568,WX10565,WX10566);
	or 	XG8228 	(WX10582,WX10579,WX10580);
	or 	XG8229 	(WX10596,WX10593,WX10594);
	or 	XG8230 	(WX10610,WX10607,WX10608);
	or 	XG8231 	(WX10624,WX10621,WX10622);
	or 	XG8232 	(WX10638,WX10635,WX10636);
	or 	XG8233 	(WX10652,WX10649,WX10650);
	or 	XG8234 	(WX10666,WX10663,WX10664);
	or 	XG8235 	(WX10680,WX10677,WX10678);
	or 	XG8236 	(WX10694,WX10691,WX10692);
	or 	XG8237 	(WX10708,WX10705,WX10706);
	or 	XG8238 	(WX10722,WX10719,WX10720);
	or 	XG8239 	(WX10736,WX10733,WX10734);
	or 	XG8240 	(WX10750,WX10747,WX10748);
	or 	XG8241 	(WX10764,WX10761,WX10762);
	or 	XG8242 	(WX10778,WX10775,WX10776);
	or 	XG8243 	(WX10792,WX10789,WX10790);
	or 	XG8244 	(WX10806,WX10803,WX10804);
	or 	XG8245 	(WX10820,WX10817,WX10818);
	nand 	XG8246 	(WX1262,II3712,II3711);
	nand 	XG8247 	(WX1261,II3705,II3704);
	nand 	XG8248 	(WX1260,II3698,II3697);
	nand 	XG8249 	(WX1259,II3691,II3690);
	nand 	XG8250 	(WX1258,II3684,II3683);
	nand 	XG8251 	(WX1257,II3677,II3676);
	nand 	XG8252 	(WX1256,II3670,II3669);
	nand 	XG8253 	(WX1255,II3663,II3662);
	nand 	XG8254 	(WX1254,II3656,II3655);
	nand 	XG8255 	(WX1253,II3649,II3648);
	nand 	XG8256 	(WX1252,II3642,II3641);
	nand 	XG8257 	(WX1251,II3635,II3634);
	nand 	XG8258 	(WX1250,II3628,II3627);
	nand 	XG8259 	(WX1249,II3621,II3620);
	nand 	XG8260 	(WX1248,II3614,II3613);
	nand 	XG8261 	(WX1247,II3607,II3606);
	nand 	XG8262 	(WX1246,II3600,II3599);
	nand 	XG8263 	(WX1245,II3593,II3592);
	nand 	XG8264 	(WX1244,II3586,II3585);
	nand 	XG8265 	(WX1243,II3579,II3578);
	nand 	XG8266 	(WX1242,II3572,II3571);
	nand 	XG8267 	(WX1241,II3565,II3564);
	nand 	XG8268 	(WX1240,II3558,II3557);
	nand 	XG8269 	(WX1239,II3551,II3550);
	nand 	XG8270 	(WX1238,II3544,II3543);
	nand 	XG8271 	(WX1237,II3537,II3536);
	nand 	XG8272 	(WX1236,II3530,II3529);
	nand 	XG8273 	(WX1235,II3523,II3522);
	nand 	XG8274 	(WX1234,II3516,II3515);
	nand 	XG8275 	(II3499,II3502,II3501);
	nand 	XG8276 	(II3484,II3487,II3486);
	nand 	XG8277 	(II3469,II3472,II3471);
	nand 	XG8278 	(WX2555,II7717,II7716);
	nand 	XG8279 	(WX2554,II7710,II7709);
	nand 	XG8280 	(WX2553,II7703,II7702);
	nand 	XG8281 	(WX2552,II7696,II7695);
	nand 	XG8282 	(WX2551,II7689,II7688);
	nand 	XG8283 	(WX2550,II7682,II7681);
	nand 	XG8284 	(WX2549,II7675,II7674);
	nand 	XG8285 	(WX2548,II7668,II7667);
	nand 	XG8286 	(WX2547,II7661,II7660);
	nand 	XG8287 	(WX2546,II7654,II7653);
	nand 	XG8288 	(WX2545,II7647,II7646);
	nand 	XG8289 	(WX2544,II7640,II7639);
	nand 	XG8290 	(WX2543,II7633,II7632);
	nand 	XG8291 	(WX2542,II7626,II7625);
	nand 	XG8292 	(WX2541,II7619,II7618);
	nand 	XG8293 	(WX2540,II7612,II7611);
	nand 	XG8294 	(WX2539,II7605,II7604);
	nand 	XG8295 	(WX2538,II7598,II7597);
	nand 	XG8296 	(WX2537,II7591,II7590);
	nand 	XG8297 	(WX2536,II7584,II7583);
	nand 	XG8298 	(WX2535,II7577,II7576);
	nand 	XG8299 	(WX2534,II7570,II7569);
	nand 	XG8300 	(WX2533,II7563,II7562);
	nand 	XG8301 	(WX2532,II7556,II7555);
	nand 	XG8302 	(WX2531,II7549,II7548);
	nand 	XG8303 	(WX2530,II7542,II7541);
	nand 	XG8304 	(WX2529,II7535,II7534);
	nand 	XG8305 	(WX2528,II7528,II7527);
	nand 	XG8306 	(WX2527,II7521,II7520);
	nand 	XG8307 	(II7504,II7507,II7506);
	nand 	XG8308 	(II7489,II7492,II7491);
	nand 	XG8309 	(II7474,II7477,II7476);
	nand 	XG8310 	(WX3848,II11722,II11721);
	nand 	XG8311 	(WX3847,II11715,II11714);
	nand 	XG8312 	(WX3846,II11708,II11707);
	nand 	XG8313 	(WX3845,II11701,II11700);
	nand 	XG8314 	(WX3844,II11694,II11693);
	nand 	XG8315 	(WX3843,II11687,II11686);
	nand 	XG8316 	(WX3842,II11680,II11679);
	nand 	XG8317 	(WX3841,II11673,II11672);
	nand 	XG8318 	(WX3840,II11666,II11665);
	nand 	XG8319 	(WX3839,II11659,II11658);
	nand 	XG8320 	(WX3838,II11652,II11651);
	nand 	XG8321 	(WX3837,II11645,II11644);
	nand 	XG8322 	(WX3836,II11638,II11637);
	nand 	XG8323 	(WX3835,II11631,II11630);
	nand 	XG8324 	(WX3834,II11624,II11623);
	nand 	XG8325 	(WX3833,II11617,II11616);
	nand 	XG8326 	(WX3832,II11610,II11609);
	nand 	XG8327 	(WX3831,II11603,II11602);
	nand 	XG8328 	(WX3830,II11596,II11595);
	nand 	XG8329 	(WX3829,II11589,II11588);
	nand 	XG8330 	(WX3828,II11582,II11581);
	nand 	XG8331 	(WX3827,II11575,II11574);
	nand 	XG8332 	(WX3826,II11568,II11567);
	nand 	XG8333 	(WX3825,II11561,II11560);
	nand 	XG8334 	(WX3824,II11554,II11553);
	nand 	XG8335 	(WX3823,II11547,II11546);
	nand 	XG8336 	(WX3822,II11540,II11539);
	nand 	XG8337 	(WX3821,II11533,II11532);
	nand 	XG8338 	(WX3820,II11526,II11525);
	nand 	XG8339 	(II11509,II11512,II11511);
	nand 	XG8340 	(II11494,II11497,II11496);
	nand 	XG8341 	(II11479,II11482,II11481);
	nand 	XG8342 	(WX5141,II15727,II15726);
	nand 	XG8343 	(WX5140,II15720,II15719);
	nand 	XG8344 	(WX5139,II15713,II15712);
	nand 	XG8345 	(WX5138,II15706,II15705);
	nand 	XG8346 	(WX5137,II15699,II15698);
	nand 	XG8347 	(WX5136,II15692,II15691);
	nand 	XG8348 	(WX5135,II15685,II15684);
	nand 	XG8349 	(WX5134,II15678,II15677);
	nand 	XG8350 	(WX5133,II15671,II15670);
	nand 	XG8351 	(WX5132,II15664,II15663);
	nand 	XG8352 	(WX5131,II15657,II15656);
	nand 	XG8353 	(WX5130,II15650,II15649);
	nand 	XG8354 	(WX5129,II15643,II15642);
	nand 	XG8355 	(WX5128,II15636,II15635);
	nand 	XG8356 	(WX5127,II15629,II15628);
	nand 	XG8357 	(WX5126,II15622,II15621);
	nand 	XG8358 	(WX5125,II15615,II15614);
	nand 	XG8359 	(WX5124,II15608,II15607);
	nand 	XG8360 	(WX5123,II15601,II15600);
	nand 	XG8361 	(WX5122,II15594,II15593);
	nand 	XG8362 	(WX5121,II15587,II15586);
	nand 	XG8363 	(WX5120,II15580,II15579);
	nand 	XG8364 	(WX5119,II15573,II15572);
	nand 	XG8365 	(WX5118,II15566,II15565);
	nand 	XG8366 	(WX5117,II15559,II15558);
	nand 	XG8367 	(WX5116,II15552,II15551);
	nand 	XG8368 	(WX5115,II15545,II15544);
	nand 	XG8369 	(WX5114,II15538,II15537);
	nand 	XG8370 	(WX5113,II15531,II15530);
	nand 	XG8371 	(II15514,II15517,II15516);
	nand 	XG8372 	(II15499,II15502,II15501);
	nand 	XG8373 	(II15484,II15487,II15486);
	nand 	XG8374 	(WX6434,II19732,II19731);
	nand 	XG8375 	(WX6433,II19725,II19724);
	nand 	XG8376 	(WX6432,II19718,II19717);
	nand 	XG8377 	(WX6431,II19711,II19710);
	nand 	XG8378 	(WX6430,II19704,II19703);
	nand 	XG8379 	(WX6429,II19697,II19696);
	nand 	XG8380 	(WX6428,II19690,II19689);
	nand 	XG8381 	(WX6427,II19683,II19682);
	nand 	XG8382 	(WX6426,II19676,II19675);
	nand 	XG8383 	(WX6425,II19669,II19668);
	nand 	XG8384 	(WX6424,II19662,II19661);
	nand 	XG8385 	(WX6423,II19655,II19654);
	nand 	XG8386 	(WX6422,II19648,II19647);
	nand 	XG8387 	(WX6421,II19641,II19640);
	nand 	XG8388 	(WX6420,II19634,II19633);
	nand 	XG8389 	(WX6419,II19627,II19626);
	nand 	XG8390 	(WX6418,II19620,II19619);
	nand 	XG8391 	(WX6417,II19613,II19612);
	nand 	XG8392 	(WX6416,II19606,II19605);
	nand 	XG8393 	(WX6415,II19599,II19598);
	nand 	XG8394 	(WX6414,II19592,II19591);
	nand 	XG8395 	(WX6413,II19585,II19584);
	nand 	XG8396 	(WX6412,II19578,II19577);
	nand 	XG8397 	(WX6411,II19571,II19570);
	nand 	XG8398 	(WX6410,II19564,II19563);
	nand 	XG8399 	(WX6409,II19557,II19556);
	nand 	XG8400 	(WX6408,II19550,II19549);
	nand 	XG8401 	(WX6407,II19543,II19542);
	nand 	XG8402 	(WX6406,II19536,II19535);
	nand 	XG8403 	(II19519,II19522,II19521);
	nand 	XG8404 	(II19504,II19507,II19506);
	nand 	XG8405 	(II19489,II19492,II19491);
	nand 	XG8406 	(WX7727,II23737,II23736);
	nand 	XG8407 	(WX7726,II23730,II23729);
	nand 	XG8408 	(WX7725,II23723,II23722);
	nand 	XG8409 	(WX7724,II23716,II23715);
	nand 	XG8410 	(WX7723,II23709,II23708);
	nand 	XG8411 	(WX7722,II23702,II23701);
	nand 	XG8412 	(WX7721,II23695,II23694);
	nand 	XG8413 	(WX7720,II23688,II23687);
	nand 	XG8414 	(WX7719,II23681,II23680);
	nand 	XG8415 	(WX7718,II23674,II23673);
	nand 	XG8416 	(WX7717,II23667,II23666);
	nand 	XG8417 	(WX7716,II23660,II23659);
	nand 	XG8418 	(WX7715,II23653,II23652);
	nand 	XG8419 	(WX7714,II23646,II23645);
	nand 	XG8420 	(WX7713,II23639,II23638);
	nand 	XG8421 	(WX7712,II23632,II23631);
	nand 	XG8422 	(WX7711,II23625,II23624);
	nand 	XG8423 	(WX7710,II23618,II23617);
	nand 	XG8424 	(WX7709,II23611,II23610);
	nand 	XG8425 	(WX7708,II23604,II23603);
	nand 	XG8426 	(WX7707,II23597,II23596);
	nand 	XG8427 	(WX7706,II23590,II23589);
	nand 	XG8428 	(WX7705,II23583,II23582);
	nand 	XG8429 	(WX7704,II23576,II23575);
	nand 	XG8430 	(WX7703,II23569,II23568);
	nand 	XG8431 	(WX7702,II23562,II23561);
	nand 	XG8432 	(WX7701,II23555,II23554);
	nand 	XG8433 	(WX7700,II23548,II23547);
	nand 	XG8434 	(WX7699,II23541,II23540);
	nand 	XG8435 	(II23524,II23527,II23526);
	nand 	XG8436 	(II23509,II23512,II23511);
	nand 	XG8437 	(II23494,II23497,II23496);
	nand 	XG8438 	(WX9020,II27742,II27741);
	nand 	XG8439 	(WX9019,II27735,II27734);
	nand 	XG8440 	(WX9018,II27728,II27727);
	nand 	XG8441 	(WX9017,II27721,II27720);
	nand 	XG8442 	(WX9016,II27714,II27713);
	nand 	XG8443 	(WX9015,II27707,II27706);
	nand 	XG8444 	(WX9014,II27700,II27699);
	nand 	XG8445 	(WX9013,II27693,II27692);
	nand 	XG8446 	(WX9012,II27686,II27685);
	nand 	XG8447 	(WX9011,II27679,II27678);
	nand 	XG8448 	(WX9010,II27672,II27671);
	nand 	XG8449 	(WX9009,II27665,II27664);
	nand 	XG8450 	(WX9008,II27658,II27657);
	nand 	XG8451 	(WX9007,II27651,II27650);
	nand 	XG8452 	(WX9006,II27644,II27643);
	nand 	XG8453 	(WX9005,II27637,II27636);
	nand 	XG8454 	(WX9004,II27630,II27629);
	nand 	XG8455 	(WX9003,II27623,II27622);
	nand 	XG8456 	(WX9002,II27616,II27615);
	nand 	XG8457 	(WX9001,II27609,II27608);
	nand 	XG8458 	(WX9000,II27602,II27601);
	nand 	XG8459 	(WX8999,II27595,II27594);
	nand 	XG8460 	(WX8998,II27588,II27587);
	nand 	XG8461 	(WX8997,II27581,II27580);
	nand 	XG8462 	(WX8996,II27574,II27573);
	nand 	XG8463 	(WX8995,II27567,II27566);
	nand 	XG8464 	(WX8994,II27560,II27559);
	nand 	XG8465 	(WX8993,II27553,II27552);
	nand 	XG8466 	(WX8992,II27546,II27545);
	nand 	XG8467 	(II27529,II27532,II27531);
	nand 	XG8468 	(II27514,II27517,II27516);
	nand 	XG8469 	(II27499,II27502,II27501);
	nand 	XG8470 	(WX10313,II31747,II31746);
	nand 	XG8471 	(WX10312,II31740,II31739);
	nand 	XG8472 	(WX10311,II31733,II31732);
	nand 	XG8473 	(WX10310,II31726,II31725);
	nand 	XG8474 	(WX10309,II31719,II31718);
	nand 	XG8475 	(WX10308,II31712,II31711);
	nand 	XG8476 	(WX10307,II31705,II31704);
	nand 	XG8477 	(WX10306,II31698,II31697);
	nand 	XG8478 	(WX10305,II31691,II31690);
	nand 	XG8479 	(WX10304,II31684,II31683);
	nand 	XG8480 	(WX10303,II31677,II31676);
	nand 	XG8481 	(WX10302,II31670,II31669);
	nand 	XG8482 	(WX10301,II31663,II31662);
	nand 	XG8483 	(WX10300,II31656,II31655);
	nand 	XG8484 	(WX10299,II31649,II31648);
	nand 	XG8485 	(WX10298,II31642,II31641);
	nand 	XG8486 	(WX10297,II31635,II31634);
	nand 	XG8487 	(WX10296,II31628,II31627);
	nand 	XG8488 	(WX10295,II31621,II31620);
	nand 	XG8489 	(WX10294,II31614,II31613);
	nand 	XG8490 	(WX10293,II31607,II31606);
	nand 	XG8491 	(WX10292,II31600,II31599);
	nand 	XG8492 	(WX10291,II31593,II31592);
	nand 	XG8493 	(WX10290,II31586,II31585);
	nand 	XG8494 	(WX10289,II31579,II31578);
	nand 	XG8495 	(WX10288,II31572,II31571);
	nand 	XG8496 	(WX10287,II31565,II31564);
	nand 	XG8497 	(WX10286,II31558,II31557);
	nand 	XG8498 	(WX10285,II31551,II31550);
	nand 	XG8499 	(II31534,II31537,II31536);
	nand 	XG8500 	(II31519,II31522,II31521);
	nand 	XG8501 	(II31504,II31507,II31506);
	nand 	XG8502 	(WX11606,II35752,II35751);
	nand 	XG8503 	(WX11605,II35745,II35744);
	nand 	XG8504 	(WX11604,II35738,II35737);
	nand 	XG8505 	(WX11603,II35731,II35730);
	nand 	XG8506 	(WX11602,II35724,II35723);
	nand 	XG8507 	(WX11601,II35717,II35716);
	nand 	XG8508 	(WX11600,II35710,II35709);
	nand 	XG8509 	(WX11599,II35703,II35702);
	nand 	XG8510 	(WX11598,II35696,II35695);
	nand 	XG8511 	(WX11597,II35689,II35688);
	nand 	XG8512 	(WX11596,II35682,II35681);
	nand 	XG8513 	(WX11595,II35675,II35674);
	nand 	XG8514 	(WX11594,II35668,II35667);
	nand 	XG8515 	(WX11593,II35661,II35660);
	nand 	XG8516 	(WX11592,II35654,II35653);
	nand 	XG8517 	(WX11591,II35647,II35646);
	nand 	XG8518 	(WX11590,II35640,II35639);
	nand 	XG8519 	(WX11589,II35633,II35632);
	nand 	XG8520 	(WX11588,II35626,II35625);
	nand 	XG8521 	(WX11587,II35619,II35618);
	nand 	XG8522 	(WX11586,II35612,II35611);
	nand 	XG8523 	(WX11585,II35605,II35604);
	nand 	XG8524 	(WX11584,II35598,II35597);
	nand 	XG8525 	(WX11583,II35591,II35590);
	nand 	XG8526 	(WX11582,II35584,II35583);
	nand 	XG8527 	(WX11581,II35577,II35576);
	nand 	XG8528 	(WX11580,II35570,II35569);
	nand 	XG8529 	(WX11579,II35563,II35562);
	nand 	XG8530 	(WX11578,II35556,II35555);
	nand 	XG8531 	(II35539,II35542,II35541);
	nand 	XG8532 	(II35524,II35527,II35526);
	nand 	XG8533 	(II35509,II35512,II35511);
	and 	XG8534 	(WX10814,WX10815,WX10820);
	and 	XG8535 	(WX10800,WX10801,WX10806);
	and 	XG8536 	(WX10786,WX10787,WX10792);
	and 	XG8537 	(WX10772,WX10773,WX10778);
	and 	XG8538 	(WX10758,WX10759,WX10764);
	and 	XG8539 	(WX10744,WX10745,WX10750);
	and 	XG8540 	(WX10730,WX10731,WX10736);
	and 	XG8541 	(WX10716,WX10717,WX10722);
	and 	XG8542 	(WX10702,WX10703,WX10708);
	and 	XG8543 	(WX10688,WX10689,WX10694);
	and 	XG8544 	(WX10674,WX10675,WX10680);
	and 	XG8545 	(WX10660,WX10661,WX10666);
	and 	XG8546 	(WX10646,WX10647,WX10652);
	and 	XG8547 	(WX10632,WX10633,WX10638);
	and 	XG8548 	(WX10618,WX10619,WX10624);
	and 	XG8549 	(WX10604,WX10605,WX10610);
	and 	XG8550 	(WX10590,WX10591,WX10596);
	and 	XG8551 	(WX10576,WX10577,WX10582);
	and 	XG8552 	(WX10562,WX10563,WX10568);
	and 	XG8553 	(WX10548,WX10549,WX10554);
	and 	XG8554 	(WX10534,WX10535,WX10540);
	and 	XG8555 	(WX10520,WX10521,WX10526);
	and 	XG8556 	(WX10506,WX10507,WX10512);
	and 	XG8557 	(WX10492,WX10493,WX10498);
	and 	XG8558 	(WX10478,WX10479,WX10484);
	and 	XG8559 	(WX10464,WX10465,WX10470);
	and 	XG8560 	(WX10450,WX10451,WX10456);
	and 	XG8561 	(WX10436,WX10437,WX10442);
	and 	XG8562 	(WX10422,WX10423,WX10428);
	and 	XG8563 	(WX10408,WX10409,WX10414);
	and 	XG8564 	(WX10394,WX10395,WX10400);
	and 	XG8565 	(WX10380,WX10381,WX10386);
	nand 	XG8566 	(II34996,II34988,WX11115);
	nand 	XG8567 	(II34965,II34957,WX11113);
	nand 	XG8568 	(II34934,II34926,WX11111);
	nand 	XG8569 	(II34903,II34895,WX11109);
	nand 	XG8570 	(II34872,II34864,WX11107);
	nand 	XG8571 	(II34841,II34833,WX11105);
	nand 	XG8572 	(II34810,II34802,WX11103);
	nand 	XG8573 	(II34779,II34771,WX11101);
	nand 	XG8574 	(II34748,II34740,WX11099);
	nand 	XG8575 	(II34717,II34709,WX11097);
	nand 	XG8576 	(II34686,II34678,WX11095);
	nand 	XG8577 	(II34655,II34647,WX11093);
	nand 	XG8578 	(II34624,II34616,WX11091);
	nand 	XG8579 	(II34593,II34585,WX11089);
	nand 	XG8580 	(II34562,II34554,WX11087);
	nand 	XG8581 	(II34531,II34523,WX11085);
	nand 	XG8582 	(II34500,II34492,WX11083);
	nand 	XG8583 	(II34469,II34461,WX11081);
	nand 	XG8584 	(II34438,II34430,WX11079);
	nand 	XG8585 	(II34407,II34399,WX11077);
	nand 	XG8586 	(II34376,II34368,WX11075);
	nand 	XG8587 	(II34345,II34337,WX11073);
	nand 	XG8588 	(II34314,II34306,WX11071);
	nand 	XG8589 	(II34283,II34275,WX11069);
	nand 	XG8590 	(II34252,II34244,WX11067);
	nand 	XG8591 	(II34221,II34213,WX11065);
	nand 	XG8592 	(II34190,II34182,WX11063);
	nand 	XG8593 	(II34159,II34151,WX11061);
	nand 	XG8594 	(II34128,II34120,WX11059);
	nand 	XG8595 	(II34097,II34089,WX11057);
	nand 	XG8596 	(II34066,II34058,WX11055);
	nand 	XG8597 	(II34035,II34027,WX11053);
	nand 	XG8598 	(II30991,II30983,WX9822);
	nand 	XG8599 	(II30960,II30952,WX9820);
	nand 	XG8600 	(II30929,II30921,WX9818);
	nand 	XG8601 	(II30898,II30890,WX9816);
	nand 	XG8602 	(II30867,II30859,WX9814);
	nand 	XG8603 	(II30836,II30828,WX9812);
	nand 	XG8604 	(II30805,II30797,WX9810);
	nand 	XG8605 	(II30774,II30766,WX9808);
	nand 	XG8606 	(II30743,II30735,WX9806);
	nand 	XG8607 	(II30712,II30704,WX9804);
	nand 	XG8608 	(II30681,II30673,WX9802);
	nand 	XG8609 	(II30650,II30642,WX9800);
	nand 	XG8610 	(II30619,II30611,WX9798);
	nand 	XG8611 	(II30588,II30580,WX9796);
	nand 	XG8612 	(II30557,II30549,WX9794);
	nand 	XG8613 	(II30526,II30518,WX9792);
	nand 	XG8614 	(II30495,II30487,WX9790);
	nand 	XG8615 	(II30464,II30456,WX9788);
	nand 	XG8616 	(II30433,II30425,WX9786);
	nand 	XG8617 	(II30402,II30394,WX9784);
	nand 	XG8618 	(II30371,II30363,WX9782);
	nand 	XG8619 	(II30340,II30332,WX9780);
	nand 	XG8620 	(II30309,II30301,WX9778);
	nand 	XG8621 	(II30278,II30270,WX9776);
	nand 	XG8622 	(II30247,II30239,WX9774);
	nand 	XG8623 	(II30216,II30208,WX9772);
	nand 	XG8624 	(II30185,II30177,WX9770);
	nand 	XG8625 	(II30154,II30146,WX9768);
	nand 	XG8626 	(II30123,II30115,WX9766);
	nand 	XG8627 	(II30092,II30084,WX9764);
	nand 	XG8628 	(II30061,II30053,WX9762);
	nand 	XG8629 	(II30030,II30022,WX9760);
	nand 	XG8630 	(II26986,II26978,WX8529);
	nand 	XG8631 	(II26955,II26947,WX8527);
	nand 	XG8632 	(II26924,II26916,WX8525);
	nand 	XG8633 	(II26893,II26885,WX8523);
	nand 	XG8634 	(II26862,II26854,WX8521);
	nand 	XG8635 	(II26831,II26823,WX8519);
	nand 	XG8636 	(II26800,II26792,WX8517);
	nand 	XG8637 	(II26769,II26761,WX8515);
	nand 	XG8638 	(II26738,II26730,WX8513);
	nand 	XG8639 	(II26707,II26699,WX8511);
	nand 	XG8640 	(II26676,II26668,WX8509);
	nand 	XG8641 	(II26645,II26637,WX8507);
	nand 	XG8642 	(II26614,II26606,WX8505);
	nand 	XG8643 	(II26583,II26575,WX8503);
	nand 	XG8644 	(II26552,II26544,WX8501);
	nand 	XG8645 	(II26521,II26513,WX8499);
	nand 	XG8646 	(II26490,II26482,WX8497);
	nand 	XG8647 	(II26459,II26451,WX8495);
	nand 	XG8648 	(II26428,II26420,WX8493);
	nand 	XG8649 	(II26397,II26389,WX8491);
	nand 	XG8650 	(II26366,II26358,WX8489);
	nand 	XG8651 	(II26335,II26327,WX8487);
	nand 	XG8652 	(II26304,II26296,WX8485);
	nand 	XG8653 	(II26273,II26265,WX8483);
	nand 	XG8654 	(II26242,II26234,WX8481);
	nand 	XG8655 	(II26211,II26203,WX8479);
	nand 	XG8656 	(II26180,II26172,WX8477);
	nand 	XG8657 	(II26149,II26141,WX8475);
	nand 	XG8658 	(II26118,II26110,WX8473);
	nand 	XG8659 	(II26087,II26079,WX8471);
	nand 	XG8660 	(II26056,II26048,WX8469);
	nand 	XG8661 	(II26025,II26017,WX8467);
	nand 	XG8662 	(II22981,II22973,WX7236);
	nand 	XG8663 	(II22950,II22942,WX7234);
	nand 	XG8664 	(II22919,II22911,WX7232);
	nand 	XG8665 	(II22888,II22880,WX7230);
	nand 	XG8666 	(II22857,II22849,WX7228);
	nand 	XG8667 	(II22826,II22818,WX7226);
	nand 	XG8668 	(II22795,II22787,WX7224);
	nand 	XG8669 	(II22764,II22756,WX7222);
	nand 	XG8670 	(II22733,II22725,WX7220);
	nand 	XG8671 	(II22702,II22694,WX7218);
	nand 	XG8672 	(II22671,II22663,WX7216);
	nand 	XG8673 	(II22640,II22632,WX7214);
	nand 	XG8674 	(II22609,II22601,WX7212);
	nand 	XG8675 	(II22578,II22570,WX7210);
	nand 	XG8676 	(II22547,II22539,WX7208);
	nand 	XG8677 	(II22516,II22508,WX7206);
	nand 	XG8678 	(II22485,II22477,WX7204);
	nand 	XG8679 	(II22454,II22446,WX7202);
	nand 	XG8680 	(II22423,II22415,WX7200);
	nand 	XG8681 	(II22392,II22384,WX7198);
	nand 	XG8682 	(II22361,II22353,WX7196);
	nand 	XG8683 	(II22330,II22322,WX7194);
	nand 	XG8684 	(II22299,II22291,WX7192);
	nand 	XG8685 	(II22268,II22260,WX7190);
	nand 	XG8686 	(II22237,II22229,WX7188);
	nand 	XG8687 	(II22206,II22198,WX7186);
	nand 	XG8688 	(II22175,II22167,WX7184);
	nand 	XG8689 	(II22144,II22136,WX7182);
	nand 	XG8690 	(II22113,II22105,WX7180);
	nand 	XG8691 	(II22082,II22074,WX7178);
	nand 	XG8692 	(II22051,II22043,WX7176);
	nand 	XG8693 	(II22020,II22012,WX7174);
	nand 	XG8694 	(II18976,II18968,WX5943);
	nand 	XG8695 	(II18945,II18937,WX5941);
	nand 	XG8696 	(II18914,II18906,WX5939);
	nand 	XG8697 	(II18883,II18875,WX5937);
	nand 	XG8698 	(II18852,II18844,WX5935);
	nand 	XG8699 	(II18821,II18813,WX5933);
	nand 	XG8700 	(II18790,II18782,WX5931);
	nand 	XG8701 	(II18759,II18751,WX5929);
	nand 	XG8702 	(II18728,II18720,WX5927);
	nand 	XG8703 	(II18697,II18689,WX5925);
	nand 	XG8704 	(II18666,II18658,WX5923);
	nand 	XG8705 	(II18635,II18627,WX5921);
	nand 	XG8706 	(II18604,II18596,WX5919);
	nand 	XG8707 	(II18573,II18565,WX5917);
	nand 	XG8708 	(II18542,II18534,WX5915);
	nand 	XG8709 	(II18511,II18503,WX5913);
	nand 	XG8710 	(II18480,II18472,WX5911);
	nand 	XG8711 	(II18449,II18441,WX5909);
	nand 	XG8712 	(II18418,II18410,WX5907);
	nand 	XG8713 	(II18387,II18379,WX5905);
	nand 	XG8714 	(II18356,II18348,WX5903);
	nand 	XG8715 	(II18325,II18317,WX5901);
	nand 	XG8716 	(II18294,II18286,WX5899);
	nand 	XG8717 	(II18263,II18255,WX5897);
	nand 	XG8718 	(II18232,II18224,WX5895);
	nand 	XG8719 	(II18201,II18193,WX5893);
	nand 	XG8720 	(II18170,II18162,WX5891);
	nand 	XG8721 	(II18139,II18131,WX5889);
	nand 	XG8722 	(II18108,II18100,WX5887);
	nand 	XG8723 	(II18077,II18069,WX5885);
	nand 	XG8724 	(II18046,II18038,WX5883);
	nand 	XG8725 	(II18015,II18007,WX5881);
	nand 	XG8726 	(II14971,II14963,WX4650);
	nand 	XG8727 	(II14940,II14932,WX4648);
	nand 	XG8728 	(II14909,II14901,WX4646);
	nand 	XG8729 	(II14878,II14870,WX4644);
	nand 	XG8730 	(II14847,II14839,WX4642);
	nand 	XG8731 	(II14816,II14808,WX4640);
	nand 	XG8732 	(II14785,II14777,WX4638);
	nand 	XG8733 	(II14754,II14746,WX4636);
	nand 	XG8734 	(II14723,II14715,WX4634);
	nand 	XG8735 	(II14692,II14684,WX4632);
	nand 	XG8736 	(II14661,II14653,WX4630);
	nand 	XG8737 	(II14630,II14622,WX4628);
	nand 	XG8738 	(II14599,II14591,WX4626);
	nand 	XG8739 	(II14568,II14560,WX4624);
	nand 	XG8740 	(II14537,II14529,WX4622);
	nand 	XG8741 	(II14506,II14498,WX4620);
	nand 	XG8742 	(II14475,II14467,WX4618);
	nand 	XG8743 	(II14444,II14436,WX4616);
	nand 	XG8744 	(II14413,II14405,WX4614);
	nand 	XG8745 	(II14382,II14374,WX4612);
	nand 	XG8746 	(II14351,II14343,WX4610);
	nand 	XG8747 	(II14320,II14312,WX4608);
	nand 	XG8748 	(II14289,II14281,WX4606);
	nand 	XG8749 	(II14258,II14250,WX4604);
	nand 	XG8750 	(II14227,II14219,WX4602);
	nand 	XG8751 	(II14196,II14188,WX4600);
	nand 	XG8752 	(II14165,II14157,WX4598);
	nand 	XG8753 	(II14134,II14126,WX4596);
	nand 	XG8754 	(II14103,II14095,WX4594);
	nand 	XG8755 	(II14072,II14064,WX4592);
	nand 	XG8756 	(II14041,II14033,WX4590);
	nand 	XG8757 	(II14010,II14002,WX4588);
	nand 	XG8758 	(II10966,II10958,WX3357);
	nand 	XG8759 	(II10935,II10927,WX3355);
	nand 	XG8760 	(II10904,II10896,WX3353);
	nand 	XG8761 	(II10873,II10865,WX3351);
	nand 	XG8762 	(II10842,II10834,WX3349);
	nand 	XG8763 	(II10811,II10803,WX3347);
	nand 	XG8764 	(II10780,II10772,WX3345);
	nand 	XG8765 	(II10749,II10741,WX3343);
	nand 	XG8766 	(II10718,II10710,WX3341);
	nand 	XG8767 	(II10687,II10679,WX3339);
	nand 	XG8768 	(II10656,II10648,WX3337);
	nand 	XG8769 	(II10625,II10617,WX3335);
	nand 	XG8770 	(II10594,II10586,WX3333);
	nand 	XG8771 	(II10563,II10555,WX3331);
	nand 	XG8772 	(II10532,II10524,WX3329);
	nand 	XG8773 	(II10501,II10493,WX3327);
	nand 	XG8774 	(II10470,II10462,WX3325);
	nand 	XG8775 	(II10439,II10431,WX3323);
	nand 	XG8776 	(II10408,II10400,WX3321);
	nand 	XG8777 	(II10377,II10369,WX3319);
	nand 	XG8778 	(II10346,II10338,WX3317);
	nand 	XG8779 	(II10315,II10307,WX3315);
	nand 	XG8780 	(II10284,II10276,WX3313);
	nand 	XG8781 	(II10253,II10245,WX3311);
	nand 	XG8782 	(II10222,II10214,WX3309);
	nand 	XG8783 	(II10191,II10183,WX3307);
	nand 	XG8784 	(II10160,II10152,WX3305);
	nand 	XG8785 	(II10129,II10121,WX3303);
	nand 	XG8786 	(II10098,II10090,WX3301);
	nand 	XG8787 	(II10067,II10059,WX3299);
	nand 	XG8788 	(II10036,II10028,WX3297);
	nand 	XG8789 	(II10005,II9997,WX3295);
	nand 	XG8790 	(II6961,II6953,WX2064);
	nand 	XG8791 	(II6930,II6922,WX2062);
	nand 	XG8792 	(II6899,II6891,WX2060);
	nand 	XG8793 	(II6868,II6860,WX2058);
	nand 	XG8794 	(II6837,II6829,WX2056);
	nand 	XG8795 	(II6806,II6798,WX2054);
	nand 	XG8796 	(II6775,II6767,WX2052);
	nand 	XG8797 	(II6744,II6736,WX2050);
	nand 	XG8798 	(II6713,II6705,WX2048);
	nand 	XG8799 	(II6682,II6674,WX2046);
	nand 	XG8800 	(II6651,II6643,WX2044);
	nand 	XG8801 	(II6620,II6612,WX2042);
	nand 	XG8802 	(II6589,II6581,WX2040);
	nand 	XG8803 	(II6558,II6550,WX2038);
	nand 	XG8804 	(II6527,II6519,WX2036);
	nand 	XG8805 	(II6496,II6488,WX2034);
	nand 	XG8806 	(II6465,II6457,WX2032);
	nand 	XG8807 	(II6434,II6426,WX2030);
	nand 	XG8808 	(II6403,II6395,WX2028);
	nand 	XG8809 	(II6372,II6364,WX2026);
	nand 	XG8810 	(II6341,II6333,WX2024);
	nand 	XG8811 	(II6310,II6302,WX2022);
	nand 	XG8812 	(II6279,II6271,WX2020);
	nand 	XG8813 	(II6248,II6240,WX2018);
	nand 	XG8814 	(II6217,II6209,WX2016);
	nand 	XG8815 	(II6186,II6178,WX2014);
	nand 	XG8816 	(II6155,II6147,WX2012);
	nand 	XG8817 	(II6124,II6116,WX2010);
	nand 	XG8818 	(II6093,II6085,WX2008);
	nand 	XG8819 	(II6062,II6054,WX2006);
	nand 	XG8820 	(II6031,II6023,WX2004);
	nand 	XG8821 	(II6000,II5992,WX2002);
	nand 	XG8822 	(II2956,II2948,WX771);
	nand 	XG8823 	(II2925,II2917,WX769);
	nand 	XG8824 	(II2894,II2886,WX767);
	nand 	XG8825 	(II2863,II2855,WX765);
	nand 	XG8826 	(II2832,II2824,WX763);
	nand 	XG8827 	(II2801,II2793,WX761);
	nand 	XG8828 	(II2770,II2762,WX759);
	nand 	XG8829 	(II2739,II2731,WX757);
	nand 	XG8830 	(II2708,II2700,WX755);
	nand 	XG8831 	(II2677,II2669,WX753);
	nand 	XG8832 	(II2646,II2638,WX751);
	nand 	XG8833 	(II2615,II2607,WX749);
	nand 	XG8834 	(II2584,II2576,WX747);
	nand 	XG8835 	(II2553,II2545,WX745);
	nand 	XG8836 	(II2522,II2514,WX743);
	nand 	XG8837 	(II2491,II2483,WX741);
	nand 	XG8838 	(II2460,II2452,WX739);
	nand 	XG8839 	(II2429,II2421,WX737);
	nand 	XG8840 	(II2398,II2390,WX735);
	nand 	XG8841 	(II2367,II2359,WX733);
	nand 	XG8842 	(II2336,II2328,WX731);
	nand 	XG8843 	(II2305,II2297,WX729);
	nand 	XG8844 	(II2274,II2266,WX727);
	nand 	XG8845 	(II2243,II2235,WX725);
	nand 	XG8846 	(II2212,II2204,WX723);
	nand 	XG8847 	(II2181,II2173,WX721);
	nand 	XG8848 	(II2150,II2142,WX719);
	nand 	XG8849 	(II2119,II2111,WX717);
	nand 	XG8850 	(II2088,II2080,WX715);
	nand 	XG8851 	(II2057,II2049,WX713);
	nand 	XG8852 	(II2026,II2018,WX711);
	nand 	XG8853 	(II1995,II1987,WX709);
	and 	XG8854 	(WX11670,WX11607,WX11579);
	and 	XG8855 	(WX11668,WX11607,WX11580);
	and 	XG8856 	(WX11666,WX11607,WX11581);
	and 	XG8857 	(WX11664,WX11607,WX11582);
	and 	XG8858 	(WX11662,WX11607,WX11583);
	and 	XG8859 	(WX11660,WX11607,WX11584);
	and 	XG8860 	(WX11658,WX11607,WX11585);
	and 	XG8861 	(WX11656,WX11607,WX11586);
	and 	XG8862 	(WX11654,WX11607,WX11587);
	and 	XG8863 	(WX11652,WX11607,WX11588);
	and 	XG8864 	(WX11650,WX11607,WX11589);
	and 	XG8865 	(WX11648,WX11607,WX11590);
	and 	XG8866 	(WX11646,WX11607,WX11591);
	and 	XG8867 	(WX11644,WX11607,WX11592);
	and 	XG8868 	(WX11642,WX11607,WX11593);
	and 	XG8869 	(WX11638,WX11607,WX11594);
	and 	XG8870 	(WX11636,WX11607,WX11595);
	and 	XG8871 	(WX11634,WX11607,WX11596);
	and 	XG8872 	(WX11632,WX11607,WX11597);
	and 	XG8873 	(WX11628,WX11607,WX11598);
	and 	XG8874 	(WX11626,WX11607,WX11599);
	and 	XG8875 	(WX11624,WX11607,WX11600);
	and 	XG8876 	(WX11622,WX11607,WX11601);
	and 	XG8877 	(WX11620,WX11607,WX11602);
	and 	XG8878 	(WX11618,WX11607,WX11603);
	and 	XG8879 	(WX11614,WX11607,WX11604);
	and 	XG8880 	(WX11612,WX11607,WX11605);
	and 	XG8881 	(WX11610,WX11607,WX11606);
	and 	XG8882 	(WX11608,WX11607,WX11578);
	and 	XG8883 	(WX10377,WX10314,WX10286);
	and 	XG8884 	(WX10375,WX10314,WX10287);
	and 	XG8885 	(WX10373,WX10314,WX10288);
	and 	XG8886 	(WX10371,WX10314,WX10289);
	and 	XG8887 	(WX10369,WX10314,WX10290);
	and 	XG8888 	(WX10367,WX10314,WX10291);
	and 	XG8889 	(WX10365,WX10314,WX10292);
	and 	XG8890 	(WX10363,WX10314,WX10293);
	and 	XG8891 	(WX10361,WX10314,WX10294);
	and 	XG8892 	(WX10359,WX10314,WX10295);
	and 	XG8893 	(WX10357,WX10314,WX10296);
	and 	XG8894 	(WX10355,WX10314,WX10297);
	and 	XG8895 	(WX10353,WX10314,WX10298);
	and 	XG8896 	(WX10351,WX10314,WX10299);
	and 	XG8897 	(WX10349,WX10314,WX10300);
	and 	XG8898 	(WX10345,WX10314,WX10301);
	and 	XG8899 	(WX10343,WX10314,WX10302);
	and 	XG8900 	(WX10341,WX10314,WX10303);
	and 	XG8901 	(WX10339,WX10314,WX10304);
	and 	XG8902 	(WX10335,WX10314,WX10305);
	and 	XG8903 	(WX10333,WX10314,WX10306);
	and 	XG8904 	(WX10331,WX10314,WX10307);
	and 	XG8905 	(WX10329,WX10314,WX10308);
	and 	XG8906 	(WX10327,WX10314,WX10309);
	and 	XG8907 	(WX10325,WX10314,WX10310);
	and 	XG8908 	(WX10321,WX10314,WX10311);
	and 	XG8909 	(WX10319,WX10314,WX10312);
	and 	XG8910 	(WX10317,WX10314,WX10313);
	and 	XG8911 	(WX10315,WX10314,WX10285);
	and 	XG8912 	(WX9084,WX9021,WX8993);
	and 	XG8913 	(WX9082,WX9021,WX8994);
	and 	XG8914 	(WX9080,WX9021,WX8995);
	and 	XG8915 	(WX9078,WX9021,WX8996);
	and 	XG8916 	(WX9076,WX9021,WX8997);
	and 	XG8917 	(WX9074,WX9021,WX8998);
	and 	XG8918 	(WX9072,WX9021,WX8999);
	and 	XG8919 	(WX9070,WX9021,WX9000);
	and 	XG8920 	(WX9068,WX9021,WX9001);
	and 	XG8921 	(WX9066,WX9021,WX9002);
	and 	XG8922 	(WX9064,WX9021,WX9003);
	and 	XG8923 	(WX9062,WX9021,WX9004);
	and 	XG8924 	(WX9060,WX9021,WX9005);
	and 	XG8925 	(WX9058,WX9021,WX9006);
	and 	XG8926 	(WX9056,WX9021,WX9007);
	and 	XG8927 	(WX9052,WX9021,WX9008);
	and 	XG8928 	(WX9050,WX9021,WX9009);
	and 	XG8929 	(WX9048,WX9021,WX9010);
	and 	XG8930 	(WX9046,WX9021,WX9011);
	and 	XG8931 	(WX9042,WX9021,WX9012);
	and 	XG8932 	(WX9040,WX9021,WX9013);
	and 	XG8933 	(WX9038,WX9021,WX9014);
	and 	XG8934 	(WX9036,WX9021,WX9015);
	and 	XG8935 	(WX9034,WX9021,WX9016);
	and 	XG8936 	(WX9032,WX9021,WX9017);
	and 	XG8937 	(WX9028,WX9021,WX9018);
	and 	XG8938 	(WX9026,WX9021,WX9019);
	and 	XG8939 	(WX9024,WX9021,WX9020);
	and 	XG8940 	(WX9022,WX9021,WX8992);
	and 	XG8941 	(WX7791,WX7728,WX7700);
	and 	XG8942 	(WX7789,WX7728,WX7701);
	and 	XG8943 	(WX7787,WX7728,WX7702);
	and 	XG8944 	(WX7785,WX7728,WX7703);
	and 	XG8945 	(WX7783,WX7728,WX7704);
	and 	XG8946 	(WX7781,WX7728,WX7705);
	and 	XG8947 	(WX7779,WX7728,WX7706);
	and 	XG8948 	(WX7777,WX7728,WX7707);
	and 	XG8949 	(WX7775,WX7728,WX7708);
	and 	XG8950 	(WX7773,WX7728,WX7709);
	and 	XG8951 	(WX7771,WX7728,WX7710);
	and 	XG8952 	(WX7769,WX7728,WX7711);
	and 	XG8953 	(WX7767,WX7728,WX7712);
	and 	XG8954 	(WX7765,WX7728,WX7713);
	and 	XG8955 	(WX7763,WX7728,WX7714);
	and 	XG8956 	(WX7759,WX7728,WX7715);
	and 	XG8957 	(WX7757,WX7728,WX7716);
	and 	XG8958 	(WX7755,WX7728,WX7717);
	and 	XG8959 	(WX7753,WX7728,WX7718);
	and 	XG8960 	(WX7749,WX7728,WX7719);
	and 	XG8961 	(WX7747,WX7728,WX7720);
	and 	XG8962 	(WX7745,WX7728,WX7721);
	and 	XG8963 	(WX7743,WX7728,WX7722);
	and 	XG8964 	(WX7741,WX7728,WX7723);
	and 	XG8965 	(WX7739,WX7728,WX7724);
	and 	XG8966 	(WX7735,WX7728,WX7725);
	and 	XG8967 	(WX7733,WX7728,WX7726);
	and 	XG8968 	(WX7731,WX7728,WX7727);
	and 	XG8969 	(WX7729,WX7728,WX7699);
	and 	XG8970 	(WX6498,WX6435,WX6407);
	and 	XG8971 	(WX6496,WX6435,WX6408);
	and 	XG8972 	(WX6494,WX6435,WX6409);
	and 	XG8973 	(WX6492,WX6435,WX6410);
	and 	XG8974 	(WX6490,WX6435,WX6411);
	and 	XG8975 	(WX6488,WX6435,WX6412);
	and 	XG8976 	(WX6486,WX6435,WX6413);
	and 	XG8977 	(WX6484,WX6435,WX6414);
	and 	XG8978 	(WX6482,WX6435,WX6415);
	and 	XG8979 	(WX6480,WX6435,WX6416);
	and 	XG8980 	(WX6478,WX6435,WX6417);
	and 	XG8981 	(WX6476,WX6435,WX6418);
	and 	XG8982 	(WX6474,WX6435,WX6419);
	and 	XG8983 	(WX6472,WX6435,WX6420);
	and 	XG8984 	(WX6470,WX6435,WX6421);
	and 	XG8985 	(WX6466,WX6435,WX6422);
	and 	XG8986 	(WX6464,WX6435,WX6423);
	and 	XG8987 	(WX6462,WX6435,WX6424);
	and 	XG8988 	(WX6460,WX6435,WX6425);
	and 	XG8989 	(WX6456,WX6435,WX6426);
	and 	XG8990 	(WX6454,WX6435,WX6427);
	and 	XG8991 	(WX6452,WX6435,WX6428);
	and 	XG8992 	(WX6450,WX6435,WX6429);
	and 	XG8993 	(WX6448,WX6435,WX6430);
	and 	XG8994 	(WX6446,WX6435,WX6431);
	and 	XG8995 	(WX6442,WX6435,WX6432);
	and 	XG8996 	(WX6440,WX6435,WX6433);
	and 	XG8997 	(WX6438,WX6435,WX6434);
	and 	XG8998 	(WX6436,WX6435,WX6406);
	and 	XG8999 	(WX5205,WX5142,WX5114);
	and 	XG9000 	(WX5203,WX5142,WX5115);
	and 	XG9001 	(WX5201,WX5142,WX5116);
	and 	XG9002 	(WX5199,WX5142,WX5117);
	and 	XG9003 	(WX5197,WX5142,WX5118);
	and 	XG9004 	(WX5195,WX5142,WX5119);
	and 	XG9005 	(WX5193,WX5142,WX5120);
	and 	XG9006 	(WX5191,WX5142,WX5121);
	and 	XG9007 	(WX5189,WX5142,WX5122);
	and 	XG9008 	(WX5187,WX5142,WX5123);
	and 	XG9009 	(WX5185,WX5142,WX5124);
	and 	XG9010 	(WX5183,WX5142,WX5125);
	and 	XG9011 	(WX5181,WX5142,WX5126);
	and 	XG9012 	(WX5179,WX5142,WX5127);
	and 	XG9013 	(WX5177,WX5142,WX5128);
	and 	XG9014 	(WX5173,WX5142,WX5129);
	and 	XG9015 	(WX5171,WX5142,WX5130);
	and 	XG9016 	(WX5169,WX5142,WX5131);
	and 	XG9017 	(WX5167,WX5142,WX5132);
	and 	XG9018 	(WX5163,WX5142,WX5133);
	and 	XG9019 	(WX5161,WX5142,WX5134);
	and 	XG9020 	(WX5159,WX5142,WX5135);
	and 	XG9021 	(WX5157,WX5142,WX5136);
	and 	XG9022 	(WX5155,WX5142,WX5137);
	and 	XG9023 	(WX5153,WX5142,WX5138);
	and 	XG9024 	(WX5149,WX5142,WX5139);
	and 	XG9025 	(WX5147,WX5142,WX5140);
	and 	XG9026 	(WX5145,WX5142,WX5141);
	and 	XG9027 	(WX5143,WX5142,WX5113);
	and 	XG9028 	(WX3912,WX3849,WX3821);
	and 	XG9029 	(WX3910,WX3849,WX3822);
	and 	XG9030 	(WX3908,WX3849,WX3823);
	and 	XG9031 	(WX3906,WX3849,WX3824);
	and 	XG9032 	(WX3904,WX3849,WX3825);
	and 	XG9033 	(WX3902,WX3849,WX3826);
	and 	XG9034 	(WX3900,WX3849,WX3827);
	and 	XG9035 	(WX3898,WX3849,WX3828);
	and 	XG9036 	(WX3896,WX3849,WX3829);
	and 	XG9037 	(WX3894,WX3849,WX3830);
	and 	XG9038 	(WX3892,WX3849,WX3831);
	and 	XG9039 	(WX3890,WX3849,WX3832);
	and 	XG9040 	(WX3888,WX3849,WX3833);
	and 	XG9041 	(WX3886,WX3849,WX3834);
	and 	XG9042 	(WX3884,WX3849,WX3835);
	and 	XG9043 	(WX3880,WX3849,WX3836);
	and 	XG9044 	(WX3878,WX3849,WX3837);
	and 	XG9045 	(WX3876,WX3849,WX3838);
	and 	XG9046 	(WX3874,WX3849,WX3839);
	and 	XG9047 	(WX3870,WX3849,WX3840);
	and 	XG9048 	(WX3868,WX3849,WX3841);
	and 	XG9049 	(WX3866,WX3849,WX3842);
	and 	XG9050 	(WX3864,WX3849,WX3843);
	and 	XG9051 	(WX3862,WX3849,WX3844);
	and 	XG9052 	(WX3860,WX3849,WX3845);
	and 	XG9053 	(WX3856,WX3849,WX3846);
	and 	XG9054 	(WX3854,WX3849,WX3847);
	and 	XG9055 	(WX3852,WX3849,WX3848);
	and 	XG9056 	(WX3850,WX3849,WX3820);
	and 	XG9057 	(WX2619,WX2556,WX2528);
	and 	XG9058 	(WX2617,WX2556,WX2529);
	and 	XG9059 	(WX2615,WX2556,WX2530);
	and 	XG9060 	(WX2613,WX2556,WX2531);
	and 	XG9061 	(WX2611,WX2556,WX2532);
	and 	XG9062 	(WX2609,WX2556,WX2533);
	and 	XG9063 	(WX2607,WX2556,WX2534);
	and 	XG9064 	(WX2605,WX2556,WX2535);
	and 	XG9065 	(WX2603,WX2556,WX2536);
	and 	XG9066 	(WX2601,WX2556,WX2537);
	and 	XG9067 	(WX2599,WX2556,WX2538);
	and 	XG9068 	(WX2597,WX2556,WX2539);
	and 	XG9069 	(WX2595,WX2556,WX2540);
	and 	XG9070 	(WX2593,WX2556,WX2541);
	and 	XG9071 	(WX2591,WX2556,WX2542);
	and 	XG9072 	(WX2587,WX2556,WX2543);
	and 	XG9073 	(WX2585,WX2556,WX2544);
	and 	XG9074 	(WX2583,WX2556,WX2545);
	and 	XG9075 	(WX2581,WX2556,WX2546);
	and 	XG9076 	(WX2577,WX2556,WX2547);
	and 	XG9077 	(WX2575,WX2556,WX2548);
	and 	XG9078 	(WX2573,WX2556,WX2549);
	and 	XG9079 	(WX2571,WX2556,WX2550);
	and 	XG9080 	(WX2569,WX2556,WX2551);
	and 	XG9081 	(WX2567,WX2556,WX2552);
	and 	XG9082 	(WX2563,WX2556,WX2553);
	and 	XG9083 	(WX2561,WX2556,WX2554);
	and 	XG9084 	(WX2559,WX2556,WX2555);
	and 	XG9085 	(WX2557,WX2556,WX2527);
	and 	XG9086 	(WX1326,WX1263,WX1235);
	and 	XG9087 	(WX1324,WX1263,WX1236);
	and 	XG9088 	(WX1322,WX1263,WX1237);
	and 	XG9089 	(WX1320,WX1263,WX1238);
	and 	XG9090 	(WX1318,WX1263,WX1239);
	and 	XG9091 	(WX1316,WX1263,WX1240);
	and 	XG9092 	(WX1314,WX1263,WX1241);
	and 	XG9093 	(WX1312,WX1263,WX1242);
	and 	XG9094 	(WX1310,WX1263,WX1243);
	and 	XG9095 	(WX1308,WX1263,WX1244);
	and 	XG9096 	(WX1306,WX1263,WX1245);
	and 	XG9097 	(WX1304,WX1263,WX1246);
	and 	XG9098 	(WX1302,WX1263,WX1247);
	and 	XG9099 	(WX1300,WX1263,WX1248);
	and 	XG9100 	(WX1298,WX1263,WX1249);
	and 	XG9101 	(WX1294,WX1263,WX1250);
	and 	XG9102 	(WX1292,WX1263,WX1251);
	and 	XG9103 	(WX1290,WX1263,WX1252);
	and 	XG9104 	(WX1288,WX1263,WX1253);
	and 	XG9105 	(WX1284,WX1263,WX1254);
	and 	XG9106 	(WX1282,WX1263,WX1255);
	and 	XG9107 	(WX1280,WX1263,WX1256);
	and 	XG9108 	(WX1278,WX1263,WX1257);
	and 	XG9109 	(WX1276,WX1263,WX1258);
	and 	XG9110 	(WX1274,WX1263,WX1259);
	and 	XG9111 	(WX1270,WX1263,WX1260);
	and 	XG9112 	(WX1268,WX1263,WX1261);
	and 	XG9113 	(WX1266,WX1263,WX1262);
	and 	XG9114 	(WX1264,WX1263,WX1234);
	nand 	XG9115 	(II3507,II3499,CRC_OUT_9_3);
	nand 	XG9116 	(II3492,II3484,CRC_OUT_9_10);
	nand 	XG9117 	(II3477,II3469,CRC_OUT_9_15);
	nand 	XG9118 	(II7512,II7504,CRC_OUT_8_3);
	nand 	XG9119 	(II7497,II7489,CRC_OUT_8_10);
	nand 	XG9120 	(II7482,II7474,CRC_OUT_8_15);
	nand 	XG9121 	(II11517,II11509,CRC_OUT_7_3);
	nand 	XG9122 	(II11502,II11494,CRC_OUT_7_10);
	nand 	XG9123 	(II11487,II11479,CRC_OUT_7_15);
	nand 	XG9124 	(II15522,II15514,CRC_OUT_6_3);
	nand 	XG9125 	(II15507,II15499,CRC_OUT_6_10);
	nand 	XG9126 	(II15492,II15484,CRC_OUT_6_15);
	nand 	XG9127 	(II19527,II19519,CRC_OUT_5_3);
	nand 	XG9128 	(II19512,II19504,CRC_OUT_5_10);
	nand 	XG9129 	(II19497,II19489,CRC_OUT_5_15);
	nand 	XG9130 	(II23532,II23524,CRC_OUT_4_3);
	nand 	XG9131 	(II23517,II23509,CRC_OUT_4_10);
	nand 	XG9132 	(II23502,II23494,CRC_OUT_4_15);
	nand 	XG9133 	(II27537,II27529,CRC_OUT_3_3);
	nand 	XG9134 	(II27522,II27514,CRC_OUT_3_10);
	nand 	XG9135 	(II27507,II27499,CRC_OUT_3_15);
	nand 	XG9136 	(II31542,II31534,CRC_OUT_2_3);
	nand 	XG9137 	(II31527,II31519,CRC_OUT_2_10);
	nand 	XG9138 	(II31512,II31504,CRC_OUT_2_15);
	nand 	XG9139 	(II35547,II35539,CRC_OUT_1_3);
	nand 	XG9140 	(II35532,II35524,CRC_OUT_1_10);
	nand 	XG9141 	(II35517,II35509,CRC_OUT_1_15);
	nand 	XG9142 	(II1997,II1995,II1987);
	nand 	XG9143 	(II2028,II2026,II2018);
	nand 	XG9144 	(II2059,II2057,II2049);
	nand 	XG9145 	(II2090,II2088,II2080);
	nand 	XG9146 	(II2121,II2119,II2111);
	nand 	XG9147 	(II2152,II2150,II2142);
	nand 	XG9148 	(II2183,II2181,II2173);
	nand 	XG9149 	(II2214,II2212,II2204);
	nand 	XG9150 	(II2245,II2243,II2235);
	nand 	XG9151 	(II2276,II2274,II2266);
	nand 	XG9152 	(II2307,II2305,II2297);
	nand 	XG9153 	(II2338,II2336,II2328);
	nand 	XG9154 	(II2369,II2367,II2359);
	nand 	XG9155 	(II2400,II2398,II2390);
	nand 	XG9156 	(II2431,II2429,II2421);
	nand 	XG9157 	(II2462,II2460,II2452);
	nand 	XG9158 	(II2493,II2491,II2483);
	nand 	XG9159 	(II2524,II2522,II2514);
	nand 	XG9160 	(II2555,II2553,II2545);
	nand 	XG9161 	(II2586,II2584,II2576);
	nand 	XG9162 	(II2617,II2615,II2607);
	nand 	XG9163 	(II2648,II2646,II2638);
	nand 	XG9164 	(II2679,II2677,II2669);
	nand 	XG9165 	(II2710,II2708,II2700);
	nand 	XG9166 	(II2741,II2739,II2731);
	nand 	XG9167 	(II2772,II2770,II2762);
	nand 	XG9168 	(II2803,II2801,II2793);
	nand 	XG9169 	(II2834,II2832,II2824);
	nand 	XG9170 	(II2865,II2863,II2855);
	nand 	XG9171 	(II2896,II2894,II2886);
	nand 	XG9172 	(II2927,II2925,II2917);
	nand 	XG9173 	(II2958,II2956,II2948);
	nand 	XG9174 	(II1996,II1995,WX709);
	nand 	XG9175 	(II2027,II2026,WX711);
	nand 	XG9176 	(II2058,II2057,WX713);
	nand 	XG9177 	(II2089,II2088,WX715);
	nand 	XG9178 	(II2120,II2119,WX717);
	nand 	XG9179 	(II2151,II2150,WX719);
	nand 	XG9180 	(II2182,II2181,WX721);
	nand 	XG9181 	(II2213,II2212,WX723);
	nand 	XG9182 	(II2244,II2243,WX725);
	nand 	XG9183 	(II2275,II2274,WX727);
	nand 	XG9184 	(II2306,II2305,WX729);
	nand 	XG9185 	(II2337,II2336,WX731);
	nand 	XG9186 	(II2368,II2367,WX733);
	nand 	XG9187 	(II2399,II2398,WX735);
	nand 	XG9188 	(II2430,II2429,WX737);
	nand 	XG9189 	(II2461,II2460,WX739);
	nand 	XG9190 	(II2492,II2491,WX741);
	nand 	XG9191 	(II2523,II2522,WX743);
	nand 	XG9192 	(II2554,II2553,WX745);
	nand 	XG9193 	(II2585,II2584,WX747);
	nand 	XG9194 	(II2616,II2615,WX749);
	nand 	XG9195 	(II2647,II2646,WX751);
	nand 	XG9196 	(II2678,II2677,WX753);
	nand 	XG9197 	(II2709,II2708,WX755);
	nand 	XG9198 	(II2740,II2739,WX757);
	nand 	XG9199 	(II2771,II2770,WX759);
	nand 	XG9200 	(II2802,II2801,WX761);
	nand 	XG9201 	(II2833,II2832,WX763);
	nand 	XG9202 	(II2864,II2863,WX765);
	nand 	XG9203 	(II2895,II2894,WX767);
	nand 	XG9204 	(II2926,II2925,WX769);
	nand 	XG9205 	(II2957,II2956,WX771);
	nand 	XG9206 	(II6002,II6000,II5992);
	nand 	XG9207 	(II6033,II6031,II6023);
	nand 	XG9208 	(II6064,II6062,II6054);
	nand 	XG9209 	(II6095,II6093,II6085);
	nand 	XG9210 	(II6126,II6124,II6116);
	nand 	XG9211 	(II6157,II6155,II6147);
	nand 	XG9212 	(II6188,II6186,II6178);
	nand 	XG9213 	(II6219,II6217,II6209);
	nand 	XG9214 	(II6250,II6248,II6240);
	nand 	XG9215 	(II6281,II6279,II6271);
	nand 	XG9216 	(II6312,II6310,II6302);
	nand 	XG9217 	(II6343,II6341,II6333);
	nand 	XG9218 	(II6374,II6372,II6364);
	nand 	XG9219 	(II6405,II6403,II6395);
	nand 	XG9220 	(II6436,II6434,II6426);
	nand 	XG9221 	(II6467,II6465,II6457);
	nand 	XG9222 	(II6498,II6496,II6488);
	nand 	XG9223 	(II6529,II6527,II6519);
	nand 	XG9224 	(II6560,II6558,II6550);
	nand 	XG9225 	(II6591,II6589,II6581);
	nand 	XG9226 	(II6622,II6620,II6612);
	nand 	XG9227 	(II6653,II6651,II6643);
	nand 	XG9228 	(II6684,II6682,II6674);
	nand 	XG9229 	(II6715,II6713,II6705);
	nand 	XG9230 	(II6746,II6744,II6736);
	nand 	XG9231 	(II6777,II6775,II6767);
	nand 	XG9232 	(II6808,II6806,II6798);
	nand 	XG9233 	(II6839,II6837,II6829);
	nand 	XG9234 	(II6870,II6868,II6860);
	nand 	XG9235 	(II6901,II6899,II6891);
	nand 	XG9236 	(II6932,II6930,II6922);
	nand 	XG9237 	(II6963,II6961,II6953);
	nand 	XG9238 	(II6001,II6000,WX2002);
	nand 	XG9239 	(II6032,II6031,WX2004);
	nand 	XG9240 	(II6063,II6062,WX2006);
	nand 	XG9241 	(II6094,II6093,WX2008);
	nand 	XG9242 	(II6125,II6124,WX2010);
	nand 	XG9243 	(II6156,II6155,WX2012);
	nand 	XG9244 	(II6187,II6186,WX2014);
	nand 	XG9245 	(II6218,II6217,WX2016);
	nand 	XG9246 	(II6249,II6248,WX2018);
	nand 	XG9247 	(II6280,II6279,WX2020);
	nand 	XG9248 	(II6311,II6310,WX2022);
	nand 	XG9249 	(II6342,II6341,WX2024);
	nand 	XG9250 	(II6373,II6372,WX2026);
	nand 	XG9251 	(II6404,II6403,WX2028);
	nand 	XG9252 	(II6435,II6434,WX2030);
	nand 	XG9253 	(II6466,II6465,WX2032);
	nand 	XG9254 	(II6497,II6496,WX2034);
	nand 	XG9255 	(II6528,II6527,WX2036);
	nand 	XG9256 	(II6559,II6558,WX2038);
	nand 	XG9257 	(II6590,II6589,WX2040);
	nand 	XG9258 	(II6621,II6620,WX2042);
	nand 	XG9259 	(II6652,II6651,WX2044);
	nand 	XG9260 	(II6683,II6682,WX2046);
	nand 	XG9261 	(II6714,II6713,WX2048);
	nand 	XG9262 	(II6745,II6744,WX2050);
	nand 	XG9263 	(II6776,II6775,WX2052);
	nand 	XG9264 	(II6807,II6806,WX2054);
	nand 	XG9265 	(II6838,II6837,WX2056);
	nand 	XG9266 	(II6869,II6868,WX2058);
	nand 	XG9267 	(II6900,II6899,WX2060);
	nand 	XG9268 	(II6931,II6930,WX2062);
	nand 	XG9269 	(II6962,II6961,WX2064);
	nand 	XG9270 	(II10007,II10005,II9997);
	nand 	XG9271 	(II10038,II10036,II10028);
	nand 	XG9272 	(II10069,II10067,II10059);
	nand 	XG9273 	(II10100,II10098,II10090);
	nand 	XG9274 	(II10131,II10129,II10121);
	nand 	XG9275 	(II10162,II10160,II10152);
	nand 	XG9276 	(II10193,II10191,II10183);
	nand 	XG9277 	(II10224,II10222,II10214);
	nand 	XG9278 	(II10255,II10253,II10245);
	nand 	XG9279 	(II10286,II10284,II10276);
	nand 	XG9280 	(II10317,II10315,II10307);
	nand 	XG9281 	(II10348,II10346,II10338);
	nand 	XG9282 	(II10379,II10377,II10369);
	nand 	XG9283 	(II10410,II10408,II10400);
	nand 	XG9284 	(II10441,II10439,II10431);
	nand 	XG9285 	(II10472,II10470,II10462);
	nand 	XG9286 	(II10503,II10501,II10493);
	nand 	XG9287 	(II10534,II10532,II10524);
	nand 	XG9288 	(II10565,II10563,II10555);
	nand 	XG9289 	(II10596,II10594,II10586);
	nand 	XG9290 	(II10627,II10625,II10617);
	nand 	XG9291 	(II10658,II10656,II10648);
	nand 	XG9292 	(II10689,II10687,II10679);
	nand 	XG9293 	(II10720,II10718,II10710);
	nand 	XG9294 	(II10751,II10749,II10741);
	nand 	XG9295 	(II10782,II10780,II10772);
	nand 	XG9296 	(II10813,II10811,II10803);
	nand 	XG9297 	(II10844,II10842,II10834);
	nand 	XG9298 	(II10875,II10873,II10865);
	nand 	XG9299 	(II10906,II10904,II10896);
	nand 	XG9300 	(II10937,II10935,II10927);
	nand 	XG9301 	(II10968,II10966,II10958);
	nand 	XG9302 	(II10006,II10005,WX3295);
	nand 	XG9303 	(II10037,II10036,WX3297);
	nand 	XG9304 	(II10068,II10067,WX3299);
	nand 	XG9305 	(II10099,II10098,WX3301);
	nand 	XG9306 	(II10130,II10129,WX3303);
	nand 	XG9307 	(II10161,II10160,WX3305);
	nand 	XG9308 	(II10192,II10191,WX3307);
	nand 	XG9309 	(II10223,II10222,WX3309);
	nand 	XG9310 	(II10254,II10253,WX3311);
	nand 	XG9311 	(II10285,II10284,WX3313);
	nand 	XG9312 	(II10316,II10315,WX3315);
	nand 	XG9313 	(II10347,II10346,WX3317);
	nand 	XG9314 	(II10378,II10377,WX3319);
	nand 	XG9315 	(II10409,II10408,WX3321);
	nand 	XG9316 	(II10440,II10439,WX3323);
	nand 	XG9317 	(II10471,II10470,WX3325);
	nand 	XG9318 	(II10502,II10501,WX3327);
	nand 	XG9319 	(II10533,II10532,WX3329);
	nand 	XG9320 	(II10564,II10563,WX3331);
	nand 	XG9321 	(II10595,II10594,WX3333);
	nand 	XG9322 	(II10626,II10625,WX3335);
	nand 	XG9323 	(II10657,II10656,WX3337);
	nand 	XG9324 	(II10688,II10687,WX3339);
	nand 	XG9325 	(II10719,II10718,WX3341);
	nand 	XG9326 	(II10750,II10749,WX3343);
	nand 	XG9327 	(II10781,II10780,WX3345);
	nand 	XG9328 	(II10812,II10811,WX3347);
	nand 	XG9329 	(II10843,II10842,WX3349);
	nand 	XG9330 	(II10874,II10873,WX3351);
	nand 	XG9331 	(II10905,II10904,WX3353);
	nand 	XG9332 	(II10936,II10935,WX3355);
	nand 	XG9333 	(II10967,II10966,WX3357);
	nand 	XG9334 	(II14012,II14010,II14002);
	nand 	XG9335 	(II14043,II14041,II14033);
	nand 	XG9336 	(II14074,II14072,II14064);
	nand 	XG9337 	(II14105,II14103,II14095);
	nand 	XG9338 	(II14136,II14134,II14126);
	nand 	XG9339 	(II14167,II14165,II14157);
	nand 	XG9340 	(II14198,II14196,II14188);
	nand 	XG9341 	(II14229,II14227,II14219);
	nand 	XG9342 	(II14260,II14258,II14250);
	nand 	XG9343 	(II14291,II14289,II14281);
	nand 	XG9344 	(II14322,II14320,II14312);
	nand 	XG9345 	(II14353,II14351,II14343);
	nand 	XG9346 	(II14384,II14382,II14374);
	nand 	XG9347 	(II14415,II14413,II14405);
	nand 	XG9348 	(II14446,II14444,II14436);
	nand 	XG9349 	(II14477,II14475,II14467);
	nand 	XG9350 	(II14508,II14506,II14498);
	nand 	XG9351 	(II14539,II14537,II14529);
	nand 	XG9352 	(II14570,II14568,II14560);
	nand 	XG9353 	(II14601,II14599,II14591);
	nand 	XG9354 	(II14632,II14630,II14622);
	nand 	XG9355 	(II14663,II14661,II14653);
	nand 	XG9356 	(II14694,II14692,II14684);
	nand 	XG9357 	(II14725,II14723,II14715);
	nand 	XG9358 	(II14756,II14754,II14746);
	nand 	XG9359 	(II14787,II14785,II14777);
	nand 	XG9360 	(II14818,II14816,II14808);
	nand 	XG9361 	(II14849,II14847,II14839);
	nand 	XG9362 	(II14880,II14878,II14870);
	nand 	XG9363 	(II14911,II14909,II14901);
	nand 	XG9364 	(II14942,II14940,II14932);
	nand 	XG9365 	(II14973,II14971,II14963);
	nand 	XG9366 	(II14011,II14010,WX4588);
	nand 	XG9367 	(II14042,II14041,WX4590);
	nand 	XG9368 	(II14073,II14072,WX4592);
	nand 	XG9369 	(II14104,II14103,WX4594);
	nand 	XG9370 	(II14135,II14134,WX4596);
	nand 	XG9371 	(II14166,II14165,WX4598);
	nand 	XG9372 	(II14197,II14196,WX4600);
	nand 	XG9373 	(II14228,II14227,WX4602);
	nand 	XG9374 	(II14259,II14258,WX4604);
	nand 	XG9375 	(II14290,II14289,WX4606);
	nand 	XG9376 	(II14321,II14320,WX4608);
	nand 	XG9377 	(II14352,II14351,WX4610);
	nand 	XG9378 	(II14383,II14382,WX4612);
	nand 	XG9379 	(II14414,II14413,WX4614);
	nand 	XG9380 	(II14445,II14444,WX4616);
	nand 	XG9381 	(II14476,II14475,WX4618);
	nand 	XG9382 	(II14507,II14506,WX4620);
	nand 	XG9383 	(II14538,II14537,WX4622);
	nand 	XG9384 	(II14569,II14568,WX4624);
	nand 	XG9385 	(II14600,II14599,WX4626);
	nand 	XG9386 	(II14631,II14630,WX4628);
	nand 	XG9387 	(II14662,II14661,WX4630);
	nand 	XG9388 	(II14693,II14692,WX4632);
	nand 	XG9389 	(II14724,II14723,WX4634);
	nand 	XG9390 	(II14755,II14754,WX4636);
	nand 	XG9391 	(II14786,II14785,WX4638);
	nand 	XG9392 	(II14817,II14816,WX4640);
	nand 	XG9393 	(II14848,II14847,WX4642);
	nand 	XG9394 	(II14879,II14878,WX4644);
	nand 	XG9395 	(II14910,II14909,WX4646);
	nand 	XG9396 	(II14941,II14940,WX4648);
	nand 	XG9397 	(II14972,II14971,WX4650);
	nand 	XG9398 	(II18017,II18015,II18007);
	nand 	XG9399 	(II18048,II18046,II18038);
	nand 	XG9400 	(II18079,II18077,II18069);
	nand 	XG9401 	(II18110,II18108,II18100);
	nand 	XG9402 	(II18141,II18139,II18131);
	nand 	XG9403 	(II18172,II18170,II18162);
	nand 	XG9404 	(II18203,II18201,II18193);
	nand 	XG9405 	(II18234,II18232,II18224);
	nand 	XG9406 	(II18265,II18263,II18255);
	nand 	XG9407 	(II18296,II18294,II18286);
	nand 	XG9408 	(II18327,II18325,II18317);
	nand 	XG9409 	(II18358,II18356,II18348);
	nand 	XG9410 	(II18389,II18387,II18379);
	nand 	XG9411 	(II18420,II18418,II18410);
	nand 	XG9412 	(II18451,II18449,II18441);
	nand 	XG9413 	(II18482,II18480,II18472);
	nand 	XG9414 	(II18513,II18511,II18503);
	nand 	XG9415 	(II18544,II18542,II18534);
	nand 	XG9416 	(II18575,II18573,II18565);
	nand 	XG9417 	(II18606,II18604,II18596);
	nand 	XG9418 	(II18637,II18635,II18627);
	nand 	XG9419 	(II18668,II18666,II18658);
	nand 	XG9420 	(II18699,II18697,II18689);
	nand 	XG9421 	(II18730,II18728,II18720);
	nand 	XG9422 	(II18761,II18759,II18751);
	nand 	XG9423 	(II18792,II18790,II18782);
	nand 	XG9424 	(II18823,II18821,II18813);
	nand 	XG9425 	(II18854,II18852,II18844);
	nand 	XG9426 	(II18885,II18883,II18875);
	nand 	XG9427 	(II18916,II18914,II18906);
	nand 	XG9428 	(II18947,II18945,II18937);
	nand 	XG9429 	(II18978,II18976,II18968);
	nand 	XG9430 	(II18016,II18015,WX5881);
	nand 	XG9431 	(II18047,II18046,WX5883);
	nand 	XG9432 	(II18078,II18077,WX5885);
	nand 	XG9433 	(II18109,II18108,WX5887);
	nand 	XG9434 	(II18140,II18139,WX5889);
	nand 	XG9435 	(II18171,II18170,WX5891);
	nand 	XG9436 	(II18202,II18201,WX5893);
	nand 	XG9437 	(II18233,II18232,WX5895);
	nand 	XG9438 	(II18264,II18263,WX5897);
	nand 	XG9439 	(II18295,II18294,WX5899);
	nand 	XG9440 	(II18326,II18325,WX5901);
	nand 	XG9441 	(II18357,II18356,WX5903);
	nand 	XG9442 	(II18388,II18387,WX5905);
	nand 	XG9443 	(II18419,II18418,WX5907);
	nand 	XG9444 	(II18450,II18449,WX5909);
	nand 	XG9445 	(II18481,II18480,WX5911);
	nand 	XG9446 	(II18512,II18511,WX5913);
	nand 	XG9447 	(II18543,II18542,WX5915);
	nand 	XG9448 	(II18574,II18573,WX5917);
	nand 	XG9449 	(II18605,II18604,WX5919);
	nand 	XG9450 	(II18636,II18635,WX5921);
	nand 	XG9451 	(II18667,II18666,WX5923);
	nand 	XG9452 	(II18698,II18697,WX5925);
	nand 	XG9453 	(II18729,II18728,WX5927);
	nand 	XG9454 	(II18760,II18759,WX5929);
	nand 	XG9455 	(II18791,II18790,WX5931);
	nand 	XG9456 	(II18822,II18821,WX5933);
	nand 	XG9457 	(II18853,II18852,WX5935);
	nand 	XG9458 	(II18884,II18883,WX5937);
	nand 	XG9459 	(II18915,II18914,WX5939);
	nand 	XG9460 	(II18946,II18945,WX5941);
	nand 	XG9461 	(II18977,II18976,WX5943);
	nand 	XG9462 	(II22022,II22020,II22012);
	nand 	XG9463 	(II22053,II22051,II22043);
	nand 	XG9464 	(II22084,II22082,II22074);
	nand 	XG9465 	(II22115,II22113,II22105);
	nand 	XG9466 	(II22146,II22144,II22136);
	nand 	XG9467 	(II22177,II22175,II22167);
	nand 	XG9468 	(II22208,II22206,II22198);
	nand 	XG9469 	(II22239,II22237,II22229);
	nand 	XG9470 	(II22270,II22268,II22260);
	nand 	XG9471 	(II22301,II22299,II22291);
	nand 	XG9472 	(II22332,II22330,II22322);
	nand 	XG9473 	(II22363,II22361,II22353);
	nand 	XG9474 	(II22394,II22392,II22384);
	nand 	XG9475 	(II22425,II22423,II22415);
	nand 	XG9476 	(II22456,II22454,II22446);
	nand 	XG9477 	(II22487,II22485,II22477);
	nand 	XG9478 	(II22518,II22516,II22508);
	nand 	XG9479 	(II22549,II22547,II22539);
	nand 	XG9480 	(II22580,II22578,II22570);
	nand 	XG9481 	(II22611,II22609,II22601);
	nand 	XG9482 	(II22642,II22640,II22632);
	nand 	XG9483 	(II22673,II22671,II22663);
	nand 	XG9484 	(II22704,II22702,II22694);
	nand 	XG9485 	(II22735,II22733,II22725);
	nand 	XG9486 	(II22766,II22764,II22756);
	nand 	XG9487 	(II22797,II22795,II22787);
	nand 	XG9488 	(II22828,II22826,II22818);
	nand 	XG9489 	(II22859,II22857,II22849);
	nand 	XG9490 	(II22890,II22888,II22880);
	nand 	XG9491 	(II22921,II22919,II22911);
	nand 	XG9492 	(II22952,II22950,II22942);
	nand 	XG9493 	(II22983,II22981,II22973);
	nand 	XG9494 	(II22021,II22020,WX7174);
	nand 	XG9495 	(II22052,II22051,WX7176);
	nand 	XG9496 	(II22083,II22082,WX7178);
	nand 	XG9497 	(II22114,II22113,WX7180);
	nand 	XG9498 	(II22145,II22144,WX7182);
	nand 	XG9499 	(II22176,II22175,WX7184);
	nand 	XG9500 	(II22207,II22206,WX7186);
	nand 	XG9501 	(II22238,II22237,WX7188);
	nand 	XG9502 	(II22269,II22268,WX7190);
	nand 	XG9503 	(II22300,II22299,WX7192);
	nand 	XG9504 	(II22331,II22330,WX7194);
	nand 	XG9505 	(II22362,II22361,WX7196);
	nand 	XG9506 	(II22393,II22392,WX7198);
	nand 	XG9507 	(II22424,II22423,WX7200);
	nand 	XG9508 	(II22455,II22454,WX7202);
	nand 	XG9509 	(II22486,II22485,WX7204);
	nand 	XG9510 	(II22517,II22516,WX7206);
	nand 	XG9511 	(II22548,II22547,WX7208);
	nand 	XG9512 	(II22579,II22578,WX7210);
	nand 	XG9513 	(II22610,II22609,WX7212);
	nand 	XG9514 	(II22641,II22640,WX7214);
	nand 	XG9515 	(II22672,II22671,WX7216);
	nand 	XG9516 	(II22703,II22702,WX7218);
	nand 	XG9517 	(II22734,II22733,WX7220);
	nand 	XG9518 	(II22765,II22764,WX7222);
	nand 	XG9519 	(II22796,II22795,WX7224);
	nand 	XG9520 	(II22827,II22826,WX7226);
	nand 	XG9521 	(II22858,II22857,WX7228);
	nand 	XG9522 	(II22889,II22888,WX7230);
	nand 	XG9523 	(II22920,II22919,WX7232);
	nand 	XG9524 	(II22951,II22950,WX7234);
	nand 	XG9525 	(II22982,II22981,WX7236);
	nand 	XG9526 	(II26027,II26025,II26017);
	nand 	XG9527 	(II26058,II26056,II26048);
	nand 	XG9528 	(II26089,II26087,II26079);
	nand 	XG9529 	(II26120,II26118,II26110);
	nand 	XG9530 	(II26151,II26149,II26141);
	nand 	XG9531 	(II26182,II26180,II26172);
	nand 	XG9532 	(II26213,II26211,II26203);
	nand 	XG9533 	(II26244,II26242,II26234);
	nand 	XG9534 	(II26275,II26273,II26265);
	nand 	XG9535 	(II26306,II26304,II26296);
	nand 	XG9536 	(II26337,II26335,II26327);
	nand 	XG9537 	(II26368,II26366,II26358);
	nand 	XG9538 	(II26399,II26397,II26389);
	nand 	XG9539 	(II26430,II26428,II26420);
	nand 	XG9540 	(II26461,II26459,II26451);
	nand 	XG9541 	(II26492,II26490,II26482);
	nand 	XG9542 	(II26523,II26521,II26513);
	nand 	XG9543 	(II26554,II26552,II26544);
	nand 	XG9544 	(II26585,II26583,II26575);
	nand 	XG9545 	(II26616,II26614,II26606);
	nand 	XG9546 	(II26647,II26645,II26637);
	nand 	XG9547 	(II26678,II26676,II26668);
	nand 	XG9548 	(II26709,II26707,II26699);
	nand 	XG9549 	(II26740,II26738,II26730);
	nand 	XG9550 	(II26771,II26769,II26761);
	nand 	XG9551 	(II26802,II26800,II26792);
	nand 	XG9552 	(II26833,II26831,II26823);
	nand 	XG9553 	(II26864,II26862,II26854);
	nand 	XG9554 	(II26895,II26893,II26885);
	nand 	XG9555 	(II26926,II26924,II26916);
	nand 	XG9556 	(II26957,II26955,II26947);
	nand 	XG9557 	(II26988,II26986,II26978);
	nand 	XG9558 	(II26026,II26025,WX8467);
	nand 	XG9559 	(II26057,II26056,WX8469);
	nand 	XG9560 	(II26088,II26087,WX8471);
	nand 	XG9561 	(II26119,II26118,WX8473);
	nand 	XG9562 	(II26150,II26149,WX8475);
	nand 	XG9563 	(II26181,II26180,WX8477);
	nand 	XG9564 	(II26212,II26211,WX8479);
	nand 	XG9565 	(II26243,II26242,WX8481);
	nand 	XG9566 	(II26274,II26273,WX8483);
	nand 	XG9567 	(II26305,II26304,WX8485);
	nand 	XG9568 	(II26336,II26335,WX8487);
	nand 	XG9569 	(II26367,II26366,WX8489);
	nand 	XG9570 	(II26398,II26397,WX8491);
	nand 	XG9571 	(II26429,II26428,WX8493);
	nand 	XG9572 	(II26460,II26459,WX8495);
	nand 	XG9573 	(II26491,II26490,WX8497);
	nand 	XG9574 	(II26522,II26521,WX8499);
	nand 	XG9575 	(II26553,II26552,WX8501);
	nand 	XG9576 	(II26584,II26583,WX8503);
	nand 	XG9577 	(II26615,II26614,WX8505);
	nand 	XG9578 	(II26646,II26645,WX8507);
	nand 	XG9579 	(II26677,II26676,WX8509);
	nand 	XG9580 	(II26708,II26707,WX8511);
	nand 	XG9581 	(II26739,II26738,WX8513);
	nand 	XG9582 	(II26770,II26769,WX8515);
	nand 	XG9583 	(II26801,II26800,WX8517);
	nand 	XG9584 	(II26832,II26831,WX8519);
	nand 	XG9585 	(II26863,II26862,WX8521);
	nand 	XG9586 	(II26894,II26893,WX8523);
	nand 	XG9587 	(II26925,II26924,WX8525);
	nand 	XG9588 	(II26956,II26955,WX8527);
	nand 	XG9589 	(II26987,II26986,WX8529);
	nand 	XG9590 	(II30032,II30030,II30022);
	nand 	XG9591 	(II30063,II30061,II30053);
	nand 	XG9592 	(II30094,II30092,II30084);
	nand 	XG9593 	(II30125,II30123,II30115);
	nand 	XG9594 	(II30156,II30154,II30146);
	nand 	XG9595 	(II30187,II30185,II30177);
	nand 	XG9596 	(II30218,II30216,II30208);
	nand 	XG9597 	(II30249,II30247,II30239);
	nand 	XG9598 	(II30280,II30278,II30270);
	nand 	XG9599 	(II30311,II30309,II30301);
	nand 	XG9600 	(II30342,II30340,II30332);
	nand 	XG9601 	(II30373,II30371,II30363);
	nand 	XG9602 	(II30404,II30402,II30394);
	nand 	XG9603 	(II30435,II30433,II30425);
	nand 	XG9604 	(II30466,II30464,II30456);
	nand 	XG9605 	(II30497,II30495,II30487);
	nand 	XG9606 	(II30528,II30526,II30518);
	nand 	XG9607 	(II30559,II30557,II30549);
	nand 	XG9608 	(II30590,II30588,II30580);
	nand 	XG9609 	(II30621,II30619,II30611);
	nand 	XG9610 	(II30652,II30650,II30642);
	nand 	XG9611 	(II30683,II30681,II30673);
	nand 	XG9612 	(II30714,II30712,II30704);
	nand 	XG9613 	(II30745,II30743,II30735);
	nand 	XG9614 	(II30776,II30774,II30766);
	nand 	XG9615 	(II30807,II30805,II30797);
	nand 	XG9616 	(II30838,II30836,II30828);
	nand 	XG9617 	(II30869,II30867,II30859);
	nand 	XG9618 	(II30900,II30898,II30890);
	nand 	XG9619 	(II30931,II30929,II30921);
	nand 	XG9620 	(II30962,II30960,II30952);
	nand 	XG9621 	(II30993,II30991,II30983);
	nand 	XG9622 	(II30031,II30030,WX9760);
	nand 	XG9623 	(II30062,II30061,WX9762);
	nand 	XG9624 	(II30093,II30092,WX9764);
	nand 	XG9625 	(II30124,II30123,WX9766);
	nand 	XG9626 	(II30155,II30154,WX9768);
	nand 	XG9627 	(II30186,II30185,WX9770);
	nand 	XG9628 	(II30217,II30216,WX9772);
	nand 	XG9629 	(II30248,II30247,WX9774);
	nand 	XG9630 	(II30279,II30278,WX9776);
	nand 	XG9631 	(II30310,II30309,WX9778);
	nand 	XG9632 	(II30341,II30340,WX9780);
	nand 	XG9633 	(II30372,II30371,WX9782);
	nand 	XG9634 	(II30403,II30402,WX9784);
	nand 	XG9635 	(II30434,II30433,WX9786);
	nand 	XG9636 	(II30465,II30464,WX9788);
	nand 	XG9637 	(II30496,II30495,WX9790);
	nand 	XG9638 	(II30527,II30526,WX9792);
	nand 	XG9639 	(II30558,II30557,WX9794);
	nand 	XG9640 	(II30589,II30588,WX9796);
	nand 	XG9641 	(II30620,II30619,WX9798);
	nand 	XG9642 	(II30651,II30650,WX9800);
	nand 	XG9643 	(II30682,II30681,WX9802);
	nand 	XG9644 	(II30713,II30712,WX9804);
	nand 	XG9645 	(II30744,II30743,WX9806);
	nand 	XG9646 	(II30775,II30774,WX9808);
	nand 	XG9647 	(II30806,II30805,WX9810);
	nand 	XG9648 	(II30837,II30836,WX9812);
	nand 	XG9649 	(II30868,II30867,WX9814);
	nand 	XG9650 	(II30899,II30898,WX9816);
	nand 	XG9651 	(II30930,II30929,WX9818);
	nand 	XG9652 	(II30961,II30960,WX9820);
	nand 	XG9653 	(II30992,II30991,WX9822);
	nand 	XG9654 	(II34037,II34035,II34027);
	nand 	XG9655 	(II34068,II34066,II34058);
	nand 	XG9656 	(II34099,II34097,II34089);
	nand 	XG9657 	(II34130,II34128,II34120);
	nand 	XG9658 	(II34161,II34159,II34151);
	nand 	XG9659 	(II34192,II34190,II34182);
	nand 	XG9660 	(II34223,II34221,II34213);
	nand 	XG9661 	(II34254,II34252,II34244);
	nand 	XG9662 	(II34285,II34283,II34275);
	nand 	XG9663 	(II34316,II34314,II34306);
	nand 	XG9664 	(II34347,II34345,II34337);
	nand 	XG9665 	(II34378,II34376,II34368);
	nand 	XG9666 	(II34409,II34407,II34399);
	nand 	XG9667 	(II34440,II34438,II34430);
	nand 	XG9668 	(II34471,II34469,II34461);
	nand 	XG9669 	(II34502,II34500,II34492);
	nand 	XG9670 	(II34533,II34531,II34523);
	nand 	XG9671 	(II34564,II34562,II34554);
	nand 	XG9672 	(II34595,II34593,II34585);
	nand 	XG9673 	(II34626,II34624,II34616);
	nand 	XG9674 	(II34657,II34655,II34647);
	nand 	XG9675 	(II34688,II34686,II34678);
	nand 	XG9676 	(II34719,II34717,II34709);
	nand 	XG9677 	(II34750,II34748,II34740);
	nand 	XG9678 	(II34781,II34779,II34771);
	nand 	XG9679 	(II34812,II34810,II34802);
	nand 	XG9680 	(II34843,II34841,II34833);
	nand 	XG9681 	(II34874,II34872,II34864);
	nand 	XG9682 	(II34905,II34903,II34895);
	nand 	XG9683 	(II34936,II34934,II34926);
	nand 	XG9684 	(II34967,II34965,II34957);
	nand 	XG9685 	(II34998,II34996,II34988);
	nand 	XG9686 	(II34036,II34035,WX11053);
	nand 	XG9687 	(II34067,II34066,WX11055);
	nand 	XG9688 	(II34098,II34097,WX11057);
	nand 	XG9689 	(II34129,II34128,WX11059);
	nand 	XG9690 	(II34160,II34159,WX11061);
	nand 	XG9691 	(II34191,II34190,WX11063);
	nand 	XG9692 	(II34222,II34221,WX11065);
	nand 	XG9693 	(II34253,II34252,WX11067);
	nand 	XG9694 	(II34284,II34283,WX11069);
	nand 	XG9695 	(II34315,II34314,WX11071);
	nand 	XG9696 	(II34346,II34345,WX11073);
	nand 	XG9697 	(II34377,II34376,WX11075);
	nand 	XG9698 	(II34408,II34407,WX11077);
	nand 	XG9699 	(II34439,II34438,WX11079);
	nand 	XG9700 	(II34470,II34469,WX11081);
	nand 	XG9701 	(II34501,II34500,WX11083);
	nand 	XG9702 	(II34532,II34531,WX11085);
	nand 	XG9703 	(II34563,II34562,WX11087);
	nand 	XG9704 	(II34594,II34593,WX11089);
	nand 	XG9705 	(II34625,II34624,WX11091);
	nand 	XG9706 	(II34656,II34655,WX11093);
	nand 	XG9707 	(II34687,II34686,WX11095);
	nand 	XG9708 	(II34718,II34717,WX11097);
	nand 	XG9709 	(II34749,II34748,WX11099);
	nand 	XG9710 	(II34780,II34779,WX11101);
	nand 	XG9711 	(II34811,II34810,WX11103);
	nand 	XG9712 	(II34842,II34841,WX11105);
	nand 	XG9713 	(II34873,II34872,WX11107);
	nand 	XG9714 	(II34904,II34903,WX11109);
	nand 	XG9715 	(II34935,II34934,WX11111);
	nand 	XG9716 	(II34966,II34965,WX11113);
	nand 	XG9717 	(II34997,II34996,WX11115);
	nand 	XG9718 	(II35519,II35517,II35509);
	nand 	XG9719 	(II35534,II35532,II35524);
	nand 	XG9720 	(II35549,II35547,II35539);
	nand 	XG9721 	(II31514,II31512,II31504);
	nand 	XG9722 	(II31529,II31527,II31519);
	nand 	XG9723 	(II31544,II31542,II31534);
	nand 	XG9724 	(II27509,II27507,II27499);
	nand 	XG9725 	(II27524,II27522,II27514);
	nand 	XG9726 	(II27539,II27537,II27529);
	nand 	XG9727 	(II23504,II23502,II23494);
	nand 	XG9728 	(II23519,II23517,II23509);
	nand 	XG9729 	(II23534,II23532,II23524);
	nand 	XG9730 	(II19499,II19497,II19489);
	nand 	XG9731 	(II19514,II19512,II19504);
	nand 	XG9732 	(II19529,II19527,II19519);
	nand 	XG9733 	(II15494,II15492,II15484);
	nand 	XG9734 	(II15509,II15507,II15499);
	nand 	XG9735 	(II15524,II15522,II15514);
	nand 	XG9736 	(II11489,II11487,II11479);
	nand 	XG9737 	(II11504,II11502,II11494);
	nand 	XG9738 	(II11519,II11517,II11509);
	nand 	XG9739 	(II7484,II7482,II7474);
	nand 	XG9740 	(II7499,II7497,II7489);
	nand 	XG9741 	(II7514,II7512,II7504);
	nand 	XG9742 	(II3479,II3477,II3469);
	nand 	XG9743 	(II3494,II3492,II3484);
	nand 	XG9744 	(II3509,II3507,II3499);
	nand 	XG9745 	(II3508,II3507,CRC_OUT_9_3);
	nand 	XG9746 	(II3493,II3492,CRC_OUT_9_10);
	nand 	XG9747 	(II3478,II3477,CRC_OUT_9_15);
	nand 	XG9748 	(II7513,II7512,CRC_OUT_8_3);
	nand 	XG9749 	(II7498,II7497,CRC_OUT_8_10);
	nand 	XG9750 	(II7483,II7482,CRC_OUT_8_15);
	nand 	XG9751 	(II11518,II11517,CRC_OUT_7_3);
	nand 	XG9752 	(II11503,II11502,CRC_OUT_7_10);
	nand 	XG9753 	(II11488,II11487,CRC_OUT_7_15);
	nand 	XG9754 	(II15523,II15522,CRC_OUT_6_3);
	nand 	XG9755 	(II15508,II15507,CRC_OUT_6_10);
	nand 	XG9756 	(II15493,II15492,CRC_OUT_6_15);
	nand 	XG9757 	(II19528,II19527,CRC_OUT_5_3);
	nand 	XG9758 	(II19513,II19512,CRC_OUT_5_10);
	nand 	XG9759 	(II19498,II19497,CRC_OUT_5_15);
	nand 	XG9760 	(II23533,II23532,CRC_OUT_4_3);
	nand 	XG9761 	(II23518,II23517,CRC_OUT_4_10);
	nand 	XG9762 	(II23503,II23502,CRC_OUT_4_15);
	nand 	XG9763 	(II27538,II27537,CRC_OUT_3_3);
	nand 	XG9764 	(II27523,II27522,CRC_OUT_3_10);
	nand 	XG9765 	(II27508,II27507,CRC_OUT_3_15);
	nand 	XG9766 	(II31543,II31542,CRC_OUT_2_3);
	nand 	XG9767 	(II31528,II31527,CRC_OUT_2_10);
	nand 	XG9768 	(II31513,II31512,CRC_OUT_2_15);
	nand 	XG9769 	(II35548,II35547,CRC_OUT_1_3);
	nand 	XG9770 	(II35533,II35532,CRC_OUT_1_10);
	nand 	XG9771 	(II35518,II35517,CRC_OUT_1_15);
	nand 	XG9772 	(II34987,II34998,II34997);
	nand 	XG9773 	(II34956,II34967,II34966);
	nand 	XG9774 	(II34925,II34936,II34935);
	nand 	XG9775 	(II34894,II34905,II34904);
	nand 	XG9776 	(II34863,II34874,II34873);
	nand 	XG9777 	(II34832,II34843,II34842);
	nand 	XG9778 	(II34801,II34812,II34811);
	nand 	XG9779 	(II34770,II34781,II34780);
	nand 	XG9780 	(II34739,II34750,II34749);
	nand 	XG9781 	(II34708,II34719,II34718);
	nand 	XG9782 	(II34677,II34688,II34687);
	nand 	XG9783 	(II34646,II34657,II34656);
	nand 	XG9784 	(II34615,II34626,II34625);
	nand 	XG9785 	(II34584,II34595,II34594);
	nand 	XG9786 	(II34553,II34564,II34563);
	nand 	XG9787 	(II34522,II34533,II34532);
	nand 	XG9788 	(II34491,II34502,II34501);
	nand 	XG9789 	(II34460,II34471,II34470);
	nand 	XG9790 	(II34429,II34440,II34439);
	nand 	XG9791 	(II34398,II34409,II34408);
	nand 	XG9792 	(II34367,II34378,II34377);
	nand 	XG9793 	(II34336,II34347,II34346);
	nand 	XG9794 	(II34305,II34316,II34315);
	nand 	XG9795 	(II34274,II34285,II34284);
	nand 	XG9796 	(II34243,II34254,II34253);
	nand 	XG9797 	(II34212,II34223,II34222);
	nand 	XG9798 	(II34181,II34192,II34191);
	nand 	XG9799 	(II34150,II34161,II34160);
	nand 	XG9800 	(II34119,II34130,II34129);
	nand 	XG9801 	(II34088,II34099,II34098);
	nand 	XG9802 	(II34057,II34068,II34067);
	nand 	XG9803 	(II34026,II34037,II34036);
	nand 	XG9804 	(II30982,II30993,II30992);
	nand 	XG9805 	(II30951,II30962,II30961);
	nand 	XG9806 	(II30920,II30931,II30930);
	nand 	XG9807 	(II30889,II30900,II30899);
	nand 	XG9808 	(II30858,II30869,II30868);
	nand 	XG9809 	(II30827,II30838,II30837);
	nand 	XG9810 	(II30796,II30807,II30806);
	nand 	XG9811 	(II30765,II30776,II30775);
	nand 	XG9812 	(II30734,II30745,II30744);
	nand 	XG9813 	(II30703,II30714,II30713);
	nand 	XG9814 	(II30672,II30683,II30682);
	nand 	XG9815 	(II30641,II30652,II30651);
	nand 	XG9816 	(II30610,II30621,II30620);
	nand 	XG9817 	(II30579,II30590,II30589);
	nand 	XG9818 	(II30548,II30559,II30558);
	nand 	XG9819 	(II30517,II30528,II30527);
	nand 	XG9820 	(II30486,II30497,II30496);
	nand 	XG9821 	(II30455,II30466,II30465);
	nand 	XG9822 	(II30424,II30435,II30434);
	nand 	XG9823 	(II30393,II30404,II30403);
	nand 	XG9824 	(II30362,II30373,II30372);
	nand 	XG9825 	(II30331,II30342,II30341);
	nand 	XG9826 	(II30300,II30311,II30310);
	nand 	XG9827 	(II30269,II30280,II30279);
	nand 	XG9828 	(II30238,II30249,II30248);
	nand 	XG9829 	(II30207,II30218,II30217);
	nand 	XG9830 	(II30176,II30187,II30186);
	nand 	XG9831 	(II30145,II30156,II30155);
	nand 	XG9832 	(II30114,II30125,II30124);
	nand 	XG9833 	(II30083,II30094,II30093);
	nand 	XG9834 	(II30052,II30063,II30062);
	nand 	XG9835 	(II30021,II30032,II30031);
	nand 	XG9836 	(II26977,II26988,II26987);
	nand 	XG9837 	(II26946,II26957,II26956);
	nand 	XG9838 	(II26915,II26926,II26925);
	nand 	XG9839 	(II26884,II26895,II26894);
	nand 	XG9840 	(II26853,II26864,II26863);
	nand 	XG9841 	(II26822,II26833,II26832);
	nand 	XG9842 	(II26791,II26802,II26801);
	nand 	XG9843 	(II26760,II26771,II26770);
	nand 	XG9844 	(II26729,II26740,II26739);
	nand 	XG9845 	(II26698,II26709,II26708);
	nand 	XG9846 	(II26667,II26678,II26677);
	nand 	XG9847 	(II26636,II26647,II26646);
	nand 	XG9848 	(II26605,II26616,II26615);
	nand 	XG9849 	(II26574,II26585,II26584);
	nand 	XG9850 	(II26543,II26554,II26553);
	nand 	XG9851 	(II26512,II26523,II26522);
	nand 	XG9852 	(II26481,II26492,II26491);
	nand 	XG9853 	(II26450,II26461,II26460);
	nand 	XG9854 	(II26419,II26430,II26429);
	nand 	XG9855 	(II26388,II26399,II26398);
	nand 	XG9856 	(II26357,II26368,II26367);
	nand 	XG9857 	(II26326,II26337,II26336);
	nand 	XG9858 	(II26295,II26306,II26305);
	nand 	XG9859 	(II26264,II26275,II26274);
	nand 	XG9860 	(II26233,II26244,II26243);
	nand 	XG9861 	(II26202,II26213,II26212);
	nand 	XG9862 	(II26171,II26182,II26181);
	nand 	XG9863 	(II26140,II26151,II26150);
	nand 	XG9864 	(II26109,II26120,II26119);
	nand 	XG9865 	(II26078,II26089,II26088);
	nand 	XG9866 	(II26047,II26058,II26057);
	nand 	XG9867 	(II26016,II26027,II26026);
	nand 	XG9868 	(II22972,II22983,II22982);
	nand 	XG9869 	(II22941,II22952,II22951);
	nand 	XG9870 	(II22910,II22921,II22920);
	nand 	XG9871 	(II22879,II22890,II22889);
	nand 	XG9872 	(II22848,II22859,II22858);
	nand 	XG9873 	(II22817,II22828,II22827);
	nand 	XG9874 	(II22786,II22797,II22796);
	nand 	XG9875 	(II22755,II22766,II22765);
	nand 	XG9876 	(II22724,II22735,II22734);
	nand 	XG9877 	(II22693,II22704,II22703);
	nand 	XG9878 	(II22662,II22673,II22672);
	nand 	XG9879 	(II22631,II22642,II22641);
	nand 	XG9880 	(II22600,II22611,II22610);
	nand 	XG9881 	(II22569,II22580,II22579);
	nand 	XG9882 	(II22538,II22549,II22548);
	nand 	XG9883 	(II22507,II22518,II22517);
	nand 	XG9884 	(II22476,II22487,II22486);
	nand 	XG9885 	(II22445,II22456,II22455);
	nand 	XG9886 	(II22414,II22425,II22424);
	nand 	XG9887 	(II22383,II22394,II22393);
	nand 	XG9888 	(II22352,II22363,II22362);
	nand 	XG9889 	(II22321,II22332,II22331);
	nand 	XG9890 	(II22290,II22301,II22300);
	nand 	XG9891 	(II22259,II22270,II22269);
	nand 	XG9892 	(II22228,II22239,II22238);
	nand 	XG9893 	(II22197,II22208,II22207);
	nand 	XG9894 	(II22166,II22177,II22176);
	nand 	XG9895 	(II22135,II22146,II22145);
	nand 	XG9896 	(II22104,II22115,II22114);
	nand 	XG9897 	(II22073,II22084,II22083);
	nand 	XG9898 	(II22042,II22053,II22052);
	nand 	XG9899 	(II22011,II22022,II22021);
	nand 	XG9900 	(II18967,II18978,II18977);
	nand 	XG9901 	(II18936,II18947,II18946);
	nand 	XG9902 	(II18905,II18916,II18915);
	nand 	XG9903 	(II18874,II18885,II18884);
	nand 	XG9904 	(II18843,II18854,II18853);
	nand 	XG9905 	(II18812,II18823,II18822);
	nand 	XG9906 	(II18781,II18792,II18791);
	nand 	XG9907 	(II18750,II18761,II18760);
	nand 	XG9908 	(II18719,II18730,II18729);
	nand 	XG9909 	(II18688,II18699,II18698);
	nand 	XG9910 	(II18657,II18668,II18667);
	nand 	XG9911 	(II18626,II18637,II18636);
	nand 	XG9912 	(II18595,II18606,II18605);
	nand 	XG9913 	(II18564,II18575,II18574);
	nand 	XG9914 	(II18533,II18544,II18543);
	nand 	XG9915 	(II18502,II18513,II18512);
	nand 	XG9916 	(II18471,II18482,II18481);
	nand 	XG9917 	(II18440,II18451,II18450);
	nand 	XG9918 	(II18409,II18420,II18419);
	nand 	XG9919 	(II18378,II18389,II18388);
	nand 	XG9920 	(II18347,II18358,II18357);
	nand 	XG9921 	(II18316,II18327,II18326);
	nand 	XG9922 	(II18285,II18296,II18295);
	nand 	XG9923 	(II18254,II18265,II18264);
	nand 	XG9924 	(II18223,II18234,II18233);
	nand 	XG9925 	(II18192,II18203,II18202);
	nand 	XG9926 	(II18161,II18172,II18171);
	nand 	XG9927 	(II18130,II18141,II18140);
	nand 	XG9928 	(II18099,II18110,II18109);
	nand 	XG9929 	(II18068,II18079,II18078);
	nand 	XG9930 	(II18037,II18048,II18047);
	nand 	XG9931 	(II18006,II18017,II18016);
	nand 	XG9932 	(II14962,II14973,II14972);
	nand 	XG9933 	(II14931,II14942,II14941);
	nand 	XG9934 	(II14900,II14911,II14910);
	nand 	XG9935 	(II14869,II14880,II14879);
	nand 	XG9936 	(II14838,II14849,II14848);
	nand 	XG9937 	(II14807,II14818,II14817);
	nand 	XG9938 	(II14776,II14787,II14786);
	nand 	XG9939 	(II14745,II14756,II14755);
	nand 	XG9940 	(II14714,II14725,II14724);
	nand 	XG9941 	(II14683,II14694,II14693);
	nand 	XG9942 	(II14652,II14663,II14662);
	nand 	XG9943 	(II14621,II14632,II14631);
	nand 	XG9944 	(II14590,II14601,II14600);
	nand 	XG9945 	(II14559,II14570,II14569);
	nand 	XG9946 	(II14528,II14539,II14538);
	nand 	XG9947 	(II14497,II14508,II14507);
	nand 	XG9948 	(II14466,II14477,II14476);
	nand 	XG9949 	(II14435,II14446,II14445);
	nand 	XG9950 	(II14404,II14415,II14414);
	nand 	XG9951 	(II14373,II14384,II14383);
	nand 	XG9952 	(II14342,II14353,II14352);
	nand 	XG9953 	(II14311,II14322,II14321);
	nand 	XG9954 	(II14280,II14291,II14290);
	nand 	XG9955 	(II14249,II14260,II14259);
	nand 	XG9956 	(II14218,II14229,II14228);
	nand 	XG9957 	(II14187,II14198,II14197);
	nand 	XG9958 	(II14156,II14167,II14166);
	nand 	XG9959 	(II14125,II14136,II14135);
	nand 	XG9960 	(II14094,II14105,II14104);
	nand 	XG9961 	(II14063,II14074,II14073);
	nand 	XG9962 	(II14032,II14043,II14042);
	nand 	XG9963 	(II14001,II14012,II14011);
	nand 	XG9964 	(II10957,II10968,II10967);
	nand 	XG9965 	(II10926,II10937,II10936);
	nand 	XG9966 	(II10895,II10906,II10905);
	nand 	XG9967 	(II10864,II10875,II10874);
	nand 	XG9968 	(II10833,II10844,II10843);
	nand 	XG9969 	(II10802,II10813,II10812);
	nand 	XG9970 	(II10771,II10782,II10781);
	nand 	XG9971 	(II10740,II10751,II10750);
	nand 	XG9972 	(II10709,II10720,II10719);
	nand 	XG9973 	(II10678,II10689,II10688);
	nand 	XG9974 	(II10647,II10658,II10657);
	nand 	XG9975 	(II10616,II10627,II10626);
	nand 	XG9976 	(II10585,II10596,II10595);
	nand 	XG9977 	(II10554,II10565,II10564);
	nand 	XG9978 	(II10523,II10534,II10533);
	nand 	XG9979 	(II10492,II10503,II10502);
	nand 	XG9980 	(II10461,II10472,II10471);
	nand 	XG9981 	(II10430,II10441,II10440);
	nand 	XG9982 	(II10399,II10410,II10409);
	nand 	XG9983 	(II10368,II10379,II10378);
	nand 	XG9984 	(II10337,II10348,II10347);
	nand 	XG9985 	(II10306,II10317,II10316);
	nand 	XG9986 	(II10275,II10286,II10285);
	nand 	XG9987 	(II10244,II10255,II10254);
	nand 	XG9988 	(II10213,II10224,II10223);
	nand 	XG9989 	(II10182,II10193,II10192);
	nand 	XG9990 	(II10151,II10162,II10161);
	nand 	XG9991 	(II10120,II10131,II10130);
	nand 	XG9992 	(II10089,II10100,II10099);
	nand 	XG9993 	(II10058,II10069,II10068);
	nand 	XG9994 	(II10027,II10038,II10037);
	nand 	XG9995 	(II9996,II10007,II10006);
	nand 	XG9996 	(II6952,II6963,II6962);
	nand 	XG9997 	(II6921,II6932,II6931);
	nand 	XG9998 	(II6890,II6901,II6900);
	nand 	XG9999 	(II6859,II6870,II6869);
	nand 	XG10000 	(II6828,II6839,II6838);
	nand 	XG10001 	(II6797,II6808,II6807);
	nand 	XG10002 	(II6766,II6777,II6776);
	nand 	XG10003 	(II6735,II6746,II6745);
	nand 	XG10004 	(II6704,II6715,II6714);
	nand 	XG10005 	(II6673,II6684,II6683);
	nand 	XG10006 	(II6642,II6653,II6652);
	nand 	XG10007 	(II6611,II6622,II6621);
	nand 	XG10008 	(II6580,II6591,II6590);
	nand 	XG10009 	(II6549,II6560,II6559);
	nand 	XG10010 	(II6518,II6529,II6528);
	nand 	XG10011 	(II6487,II6498,II6497);
	nand 	XG10012 	(II6456,II6467,II6466);
	nand 	XG10013 	(II6425,II6436,II6435);
	nand 	XG10014 	(II6394,II6405,II6404);
	nand 	XG10015 	(II6363,II6374,II6373);
	nand 	XG10016 	(II6332,II6343,II6342);
	nand 	XG10017 	(II6301,II6312,II6311);
	nand 	XG10018 	(II6270,II6281,II6280);
	nand 	XG10019 	(II6239,II6250,II6249);
	nand 	XG10020 	(II6208,II6219,II6218);
	nand 	XG10021 	(II6177,II6188,II6187);
	nand 	XG10022 	(II6146,II6157,II6156);
	nand 	XG10023 	(II6115,II6126,II6125);
	nand 	XG10024 	(II6084,II6095,II6094);
	nand 	XG10025 	(II6053,II6064,II6063);
	nand 	XG10026 	(II6022,II6033,II6032);
	nand 	XG10027 	(II5991,II6002,II6001);
	nand 	XG10028 	(II2947,II2958,II2957);
	nand 	XG10029 	(II2916,II2927,II2926);
	nand 	XG10030 	(II2885,II2896,II2895);
	nand 	XG10031 	(II2854,II2865,II2864);
	nand 	XG10032 	(II2823,II2834,II2833);
	nand 	XG10033 	(II2792,II2803,II2802);
	nand 	XG10034 	(II2761,II2772,II2771);
	nand 	XG10035 	(II2730,II2741,II2740);
	nand 	XG10036 	(II2699,II2710,II2709);
	nand 	XG10037 	(II2668,II2679,II2678);
	nand 	XG10038 	(II2637,II2648,II2647);
	nand 	XG10039 	(II2606,II2617,II2616);
	nand 	XG10040 	(II2575,II2586,II2585);
	nand 	XG10041 	(II2544,II2555,II2554);
	nand 	XG10042 	(II2513,II2524,II2523);
	nand 	XG10043 	(II2482,II2493,II2492);
	nand 	XG10044 	(II2451,II2462,II2461);
	nand 	XG10045 	(II2420,II2431,II2430);
	nand 	XG10046 	(II2389,II2400,II2399);
	nand 	XG10047 	(II2358,II2369,II2368);
	nand 	XG10048 	(II2327,II2338,II2337);
	nand 	XG10049 	(II2296,II2307,II2306);
	nand 	XG10050 	(II2265,II2276,II2275);
	nand 	XG10051 	(II2234,II2245,II2244);
	nand 	XG10052 	(II2203,II2214,II2213);
	nand 	XG10053 	(II2172,II2183,II2182);
	nand 	XG10054 	(II2141,II2152,II2151);
	nand 	XG10055 	(II2110,II2121,II2120);
	nand 	XG10056 	(II2079,II2090,II2089);
	nand 	XG10057 	(II2048,II2059,II2058);
	nand 	XG10058 	(II2017,II2028,II2027);
	nand 	XG10059 	(II1986,II1997,II1996);
	nand 	XG10060 	(WX1233,II3509,II3508);
	nand 	XG10061 	(WX1232,II3494,II3493);
	nand 	XG10062 	(WX1231,II3479,II3478);
	nand 	XG10063 	(WX2526,II7514,II7513);
	nand 	XG10064 	(WX2525,II7499,II7498);
	nand 	XG10065 	(WX2524,II7484,II7483);
	nand 	XG10066 	(WX3819,II11519,II11518);
	nand 	XG10067 	(WX3818,II11504,II11503);
	nand 	XG10068 	(WX3817,II11489,II11488);
	nand 	XG10069 	(WX5112,II15524,II15523);
	nand 	XG10070 	(WX5111,II15509,II15508);
	nand 	XG10071 	(WX5110,II15494,II15493);
	nand 	XG10072 	(WX6405,II19529,II19528);
	nand 	XG10073 	(WX6404,II19514,II19513);
	nand 	XG10074 	(WX6403,II19499,II19498);
	nand 	XG10075 	(WX7698,II23534,II23533);
	nand 	XG10076 	(WX7697,II23519,II23518);
	nand 	XG10077 	(WX7696,II23504,II23503);
	nand 	XG10078 	(WX8991,II27539,II27538);
	nand 	XG10079 	(WX8990,II27524,II27523);
	nand 	XG10080 	(WX8989,II27509,II27508);
	nand 	XG10081 	(WX10284,II31544,II31543);
	nand 	XG10082 	(WX10283,II31529,II31528);
	nand 	XG10083 	(WX10282,II31514,II31513);
	nand 	XG10084 	(WX11577,II35549,II35548);
	nand 	XG10085 	(WX11576,II35534,II35533);
	nand 	XG10086 	(WX11575,II35519,II35518);
	nand 	XG10087 	(II35011,II35003,II34987);
	nand 	XG10088 	(II34980,II34972,II34956);
	nand 	XG10089 	(II34949,II34941,II34925);
	nand 	XG10090 	(II34918,II34910,II34894);
	nand 	XG10091 	(II34887,II34879,II34863);
	nand 	XG10092 	(II34856,II34848,II34832);
	nand 	XG10093 	(II34825,II34817,II34801);
	nand 	XG10094 	(II34794,II34786,II34770);
	nand 	XG10095 	(II34763,II34755,II34739);
	nand 	XG10096 	(II34732,II34724,II34708);
	nand 	XG10097 	(II34701,II34693,II34677);
	nand 	XG10098 	(II34670,II34662,II34646);
	nand 	XG10099 	(II34639,II34631,II34615);
	nand 	XG10100 	(II34608,II34600,II34584);
	nand 	XG10101 	(II34577,II34569,II34553);
	nand 	XG10102 	(II34546,II34538,II34522);
	nand 	XG10103 	(II34515,II34507,II34491);
	nand 	XG10104 	(II34484,II34476,II34460);
	nand 	XG10105 	(II34453,II34445,II34429);
	nand 	XG10106 	(II34422,II34414,II34398);
	nand 	XG10107 	(II34391,II34383,II34367);
	nand 	XG10108 	(II34360,II34352,II34336);
	nand 	XG10109 	(II34329,II34321,II34305);
	nand 	XG10110 	(II34298,II34290,II34274);
	nand 	XG10111 	(II34267,II34259,II34243);
	nand 	XG10112 	(II34236,II34228,II34212);
	nand 	XG10113 	(II34205,II34197,II34181);
	nand 	XG10114 	(II34174,II34166,II34150);
	nand 	XG10115 	(II34143,II34135,II34119);
	nand 	XG10116 	(II34112,II34104,II34088);
	nand 	XG10117 	(II34081,II34073,II34057);
	nand 	XG10118 	(II34050,II34042,II34026);
	nand 	XG10119 	(II31006,II30998,II30982);
	nand 	XG10120 	(II30975,II30967,II30951);
	nand 	XG10121 	(II30944,II30936,II30920);
	nand 	XG10122 	(II30913,II30905,II30889);
	nand 	XG10123 	(II30882,II30874,II30858);
	nand 	XG10124 	(II30851,II30843,II30827);
	nand 	XG10125 	(II30820,II30812,II30796);
	nand 	XG10126 	(II30789,II30781,II30765);
	nand 	XG10127 	(II30758,II30750,II30734);
	nand 	XG10128 	(II30727,II30719,II30703);
	nand 	XG10129 	(II30696,II30688,II30672);
	nand 	XG10130 	(II30665,II30657,II30641);
	nand 	XG10131 	(II30634,II30626,II30610);
	nand 	XG10132 	(II30603,II30595,II30579);
	nand 	XG10133 	(II30572,II30564,II30548);
	nand 	XG10134 	(II30541,II30533,II30517);
	nand 	XG10135 	(II30510,II30502,II30486);
	nand 	XG10136 	(II30479,II30471,II30455);
	nand 	XG10137 	(II30448,II30440,II30424);
	nand 	XG10138 	(II30417,II30409,II30393);
	nand 	XG10139 	(II30386,II30378,II30362);
	nand 	XG10140 	(II30355,II30347,II30331);
	nand 	XG10141 	(II30324,II30316,II30300);
	nand 	XG10142 	(II30293,II30285,II30269);
	nand 	XG10143 	(II30262,II30254,II30238);
	nand 	XG10144 	(II30231,II30223,II30207);
	nand 	XG10145 	(II30200,II30192,II30176);
	nand 	XG10146 	(II30169,II30161,II30145);
	nand 	XG10147 	(II30138,II30130,II30114);
	nand 	XG10148 	(II30107,II30099,II30083);
	nand 	XG10149 	(II30076,II30068,II30052);
	nand 	XG10150 	(II30045,II30037,II30021);
	nand 	XG10151 	(II27001,II26993,II26977);
	nand 	XG10152 	(II26970,II26962,II26946);
	nand 	XG10153 	(II26939,II26931,II26915);
	nand 	XG10154 	(II26908,II26900,II26884);
	nand 	XG10155 	(II26877,II26869,II26853);
	nand 	XG10156 	(II26846,II26838,II26822);
	nand 	XG10157 	(II26815,II26807,II26791);
	nand 	XG10158 	(II26784,II26776,II26760);
	nand 	XG10159 	(II26753,II26745,II26729);
	nand 	XG10160 	(II26722,II26714,II26698);
	nand 	XG10161 	(II26691,II26683,II26667);
	nand 	XG10162 	(II26660,II26652,II26636);
	nand 	XG10163 	(II26629,II26621,II26605);
	nand 	XG10164 	(II26598,II26590,II26574);
	nand 	XG10165 	(II26567,II26559,II26543);
	nand 	XG10166 	(II26536,II26528,II26512);
	nand 	XG10167 	(II26505,II26497,II26481);
	nand 	XG10168 	(II26474,II26466,II26450);
	nand 	XG10169 	(II26443,II26435,II26419);
	nand 	XG10170 	(II26412,II26404,II26388);
	nand 	XG10171 	(II26381,II26373,II26357);
	nand 	XG10172 	(II26350,II26342,II26326);
	nand 	XG10173 	(II26319,II26311,II26295);
	nand 	XG10174 	(II26288,II26280,II26264);
	nand 	XG10175 	(II26257,II26249,II26233);
	nand 	XG10176 	(II26226,II26218,II26202);
	nand 	XG10177 	(II26195,II26187,II26171);
	nand 	XG10178 	(II26164,II26156,II26140);
	nand 	XG10179 	(II26133,II26125,II26109);
	nand 	XG10180 	(II26102,II26094,II26078);
	nand 	XG10181 	(II26071,II26063,II26047);
	nand 	XG10182 	(II26040,II26032,II26016);
	nand 	XG10183 	(II22996,II22988,II22972);
	nand 	XG10184 	(II22965,II22957,II22941);
	nand 	XG10185 	(II22934,II22926,II22910);
	nand 	XG10186 	(II22903,II22895,II22879);
	nand 	XG10187 	(II22872,II22864,II22848);
	nand 	XG10188 	(II22841,II22833,II22817);
	nand 	XG10189 	(II22810,II22802,II22786);
	nand 	XG10190 	(II22779,II22771,II22755);
	nand 	XG10191 	(II22748,II22740,II22724);
	nand 	XG10192 	(II22717,II22709,II22693);
	nand 	XG10193 	(II22686,II22678,II22662);
	nand 	XG10194 	(II22655,II22647,II22631);
	nand 	XG10195 	(II22624,II22616,II22600);
	nand 	XG10196 	(II22593,II22585,II22569);
	nand 	XG10197 	(II22562,II22554,II22538);
	nand 	XG10198 	(II22531,II22523,II22507);
	nand 	XG10199 	(II22500,II22492,II22476);
	nand 	XG10200 	(II22469,II22461,II22445);
	nand 	XG10201 	(II22438,II22430,II22414);
	nand 	XG10202 	(II22407,II22399,II22383);
	nand 	XG10203 	(II22376,II22368,II22352);
	nand 	XG10204 	(II22345,II22337,II22321);
	nand 	XG10205 	(II22314,II22306,II22290);
	nand 	XG10206 	(II22283,II22275,II22259);
	nand 	XG10207 	(II22252,II22244,II22228);
	nand 	XG10208 	(II22221,II22213,II22197);
	nand 	XG10209 	(II22190,II22182,II22166);
	nand 	XG10210 	(II22159,II22151,II22135);
	nand 	XG10211 	(II22128,II22120,II22104);
	nand 	XG10212 	(II22097,II22089,II22073);
	nand 	XG10213 	(II22066,II22058,II22042);
	nand 	XG10214 	(II22035,II22027,II22011);
	nand 	XG10215 	(II18991,II18983,II18967);
	nand 	XG10216 	(II18960,II18952,II18936);
	nand 	XG10217 	(II18929,II18921,II18905);
	nand 	XG10218 	(II18898,II18890,II18874);
	nand 	XG10219 	(II18867,II18859,II18843);
	nand 	XG10220 	(II18836,II18828,II18812);
	nand 	XG10221 	(II18805,II18797,II18781);
	nand 	XG10222 	(II18774,II18766,II18750);
	nand 	XG10223 	(II18743,II18735,II18719);
	nand 	XG10224 	(II18712,II18704,II18688);
	nand 	XG10225 	(II18681,II18673,II18657);
	nand 	XG10226 	(II18650,II18642,II18626);
	nand 	XG10227 	(II18619,II18611,II18595);
	nand 	XG10228 	(II18588,II18580,II18564);
	nand 	XG10229 	(II18557,II18549,II18533);
	nand 	XG10230 	(II18526,II18518,II18502);
	nand 	XG10231 	(II18495,II18487,II18471);
	nand 	XG10232 	(II18464,II18456,II18440);
	nand 	XG10233 	(II18433,II18425,II18409);
	nand 	XG10234 	(II18402,II18394,II18378);
	nand 	XG10235 	(II18371,II18363,II18347);
	nand 	XG10236 	(II18340,II18332,II18316);
	nand 	XG10237 	(II18309,II18301,II18285);
	nand 	XG10238 	(II18278,II18270,II18254);
	nand 	XG10239 	(II18247,II18239,II18223);
	nand 	XG10240 	(II18216,II18208,II18192);
	nand 	XG10241 	(II18185,II18177,II18161);
	nand 	XG10242 	(II18154,II18146,II18130);
	nand 	XG10243 	(II18123,II18115,II18099);
	nand 	XG10244 	(II18092,II18084,II18068);
	nand 	XG10245 	(II18061,II18053,II18037);
	nand 	XG10246 	(II18030,II18022,II18006);
	nand 	XG10247 	(II14986,II14978,II14962);
	nand 	XG10248 	(II14955,II14947,II14931);
	nand 	XG10249 	(II14924,II14916,II14900);
	nand 	XG10250 	(II14893,II14885,II14869);
	nand 	XG10251 	(II14862,II14854,II14838);
	nand 	XG10252 	(II14831,II14823,II14807);
	nand 	XG10253 	(II14800,II14792,II14776);
	nand 	XG10254 	(II14769,II14761,II14745);
	nand 	XG10255 	(II14738,II14730,II14714);
	nand 	XG10256 	(II14707,II14699,II14683);
	nand 	XG10257 	(II14676,II14668,II14652);
	nand 	XG10258 	(II14645,II14637,II14621);
	nand 	XG10259 	(II14614,II14606,II14590);
	nand 	XG10260 	(II14583,II14575,II14559);
	nand 	XG10261 	(II14552,II14544,II14528);
	nand 	XG10262 	(II14521,II14513,II14497);
	nand 	XG10263 	(II14490,II14482,II14466);
	nand 	XG10264 	(II14459,II14451,II14435);
	nand 	XG10265 	(II14428,II14420,II14404);
	nand 	XG10266 	(II14397,II14389,II14373);
	nand 	XG10267 	(II14366,II14358,II14342);
	nand 	XG10268 	(II14335,II14327,II14311);
	nand 	XG10269 	(II14304,II14296,II14280);
	nand 	XG10270 	(II14273,II14265,II14249);
	nand 	XG10271 	(II14242,II14234,II14218);
	nand 	XG10272 	(II14211,II14203,II14187);
	nand 	XG10273 	(II14180,II14172,II14156);
	nand 	XG10274 	(II14149,II14141,II14125);
	nand 	XG10275 	(II14118,II14110,II14094);
	nand 	XG10276 	(II14087,II14079,II14063);
	nand 	XG10277 	(II14056,II14048,II14032);
	nand 	XG10278 	(II14025,II14017,II14001);
	nand 	XG10279 	(II10981,II10973,II10957);
	nand 	XG10280 	(II10950,II10942,II10926);
	nand 	XG10281 	(II10919,II10911,II10895);
	nand 	XG10282 	(II10888,II10880,II10864);
	nand 	XG10283 	(II10857,II10849,II10833);
	nand 	XG10284 	(II10826,II10818,II10802);
	nand 	XG10285 	(II10795,II10787,II10771);
	nand 	XG10286 	(II10764,II10756,II10740);
	nand 	XG10287 	(II10733,II10725,II10709);
	nand 	XG10288 	(II10702,II10694,II10678);
	nand 	XG10289 	(II10671,II10663,II10647);
	nand 	XG10290 	(II10640,II10632,II10616);
	nand 	XG10291 	(II10609,II10601,II10585);
	nand 	XG10292 	(II10578,II10570,II10554);
	nand 	XG10293 	(II10547,II10539,II10523);
	nand 	XG10294 	(II10516,II10508,II10492);
	nand 	XG10295 	(II10485,II10477,II10461);
	nand 	XG10296 	(II10454,II10446,II10430);
	nand 	XG10297 	(II10423,II10415,II10399);
	nand 	XG10298 	(II10392,II10384,II10368);
	nand 	XG10299 	(II10361,II10353,II10337);
	nand 	XG10300 	(II10330,II10322,II10306);
	nand 	XG10301 	(II10299,II10291,II10275);
	nand 	XG10302 	(II10268,II10260,II10244);
	nand 	XG10303 	(II10237,II10229,II10213);
	nand 	XG10304 	(II10206,II10198,II10182);
	nand 	XG10305 	(II10175,II10167,II10151);
	nand 	XG10306 	(II10144,II10136,II10120);
	nand 	XG10307 	(II10113,II10105,II10089);
	nand 	XG10308 	(II10082,II10074,II10058);
	nand 	XG10309 	(II10051,II10043,II10027);
	nand 	XG10310 	(II10020,II10012,II9996);
	nand 	XG10311 	(II6976,II6968,II6952);
	nand 	XG10312 	(II6945,II6937,II6921);
	nand 	XG10313 	(II6914,II6906,II6890);
	nand 	XG10314 	(II6883,II6875,II6859);
	nand 	XG10315 	(II6852,II6844,II6828);
	nand 	XG10316 	(II6821,II6813,II6797);
	nand 	XG10317 	(II6790,II6782,II6766);
	nand 	XG10318 	(II6759,II6751,II6735);
	nand 	XG10319 	(II6728,II6720,II6704);
	nand 	XG10320 	(II6697,II6689,II6673);
	nand 	XG10321 	(II6666,II6658,II6642);
	nand 	XG10322 	(II6635,II6627,II6611);
	nand 	XG10323 	(II6604,II6596,II6580);
	nand 	XG10324 	(II6573,II6565,II6549);
	nand 	XG10325 	(II6542,II6534,II6518);
	nand 	XG10326 	(II6511,II6503,II6487);
	nand 	XG10327 	(II6480,II6472,II6456);
	nand 	XG10328 	(II6449,II6441,II6425);
	nand 	XG10329 	(II6418,II6410,II6394);
	nand 	XG10330 	(II6387,II6379,II6363);
	nand 	XG10331 	(II6356,II6348,II6332);
	nand 	XG10332 	(II6325,II6317,II6301);
	nand 	XG10333 	(II6294,II6286,II6270);
	nand 	XG10334 	(II6263,II6255,II6239);
	nand 	XG10335 	(II6232,II6224,II6208);
	nand 	XG10336 	(II6201,II6193,II6177);
	nand 	XG10337 	(II6170,II6162,II6146);
	nand 	XG10338 	(II6139,II6131,II6115);
	nand 	XG10339 	(II6108,II6100,II6084);
	nand 	XG10340 	(II6077,II6069,II6053);
	nand 	XG10341 	(II6046,II6038,II6022);
	nand 	XG10342 	(II6015,II6007,II5991);
	nand 	XG10343 	(II2971,II2963,II2947);
	nand 	XG10344 	(II2940,II2932,II2916);
	nand 	XG10345 	(II2909,II2901,II2885);
	nand 	XG10346 	(II2878,II2870,II2854);
	nand 	XG10347 	(II2847,II2839,II2823);
	nand 	XG10348 	(II2816,II2808,II2792);
	nand 	XG10349 	(II2785,II2777,II2761);
	nand 	XG10350 	(II2754,II2746,II2730);
	nand 	XG10351 	(II2723,II2715,II2699);
	nand 	XG10352 	(II2692,II2684,II2668);
	nand 	XG10353 	(II2661,II2653,II2637);
	nand 	XG10354 	(II2630,II2622,II2606);
	nand 	XG10355 	(II2599,II2591,II2575);
	nand 	XG10356 	(II2568,II2560,II2544);
	nand 	XG10357 	(II2537,II2529,II2513);
	nand 	XG10358 	(II2506,II2498,II2482);
	nand 	XG10359 	(II2475,II2467,II2451);
	nand 	XG10360 	(II2444,II2436,II2420);
	nand 	XG10361 	(II2413,II2405,II2389);
	nand 	XG10362 	(II2382,II2374,II2358);
	nand 	XG10363 	(II2351,II2343,II2327);
	nand 	XG10364 	(II2320,II2312,II2296);
	nand 	XG10365 	(II2289,II2281,II2265);
	nand 	XG10366 	(II2258,II2250,II2234);
	nand 	XG10367 	(II2227,II2219,II2203);
	nand 	XG10368 	(II2196,II2188,II2172);
	nand 	XG10369 	(II2165,II2157,II2141);
	nand 	XG10370 	(II2134,II2126,II2110);
	nand 	XG10371 	(II2103,II2095,II2079);
	nand 	XG10372 	(II2072,II2064,II2048);
	nand 	XG10373 	(II2041,II2033,II2017);
	nand 	XG10374 	(II2010,II2002,II1986);
	and 	XG10375 	(WX11640,WX11607,WX11575);
	and 	XG10376 	(WX11630,WX11607,WX11576);
	and 	XG10377 	(WX11616,WX11607,WX11577);
	and 	XG10378 	(WX10347,WX10314,WX10282);
	and 	XG10379 	(WX10337,WX10314,WX10283);
	and 	XG10380 	(WX10323,WX10314,WX10284);
	and 	XG10381 	(WX9054,WX9021,WX8989);
	and 	XG10382 	(WX9044,WX9021,WX8990);
	and 	XG10383 	(WX9030,WX9021,WX8991);
	and 	XG10384 	(WX7761,WX7728,WX7696);
	and 	XG10385 	(WX7751,WX7728,WX7697);
	and 	XG10386 	(WX7737,WX7728,WX7698);
	and 	XG10387 	(WX6468,WX6435,WX6403);
	and 	XG10388 	(WX6458,WX6435,WX6404);
	and 	XG10389 	(WX6444,WX6435,WX6405);
	and 	XG10390 	(WX5175,WX5142,WX5110);
	and 	XG10391 	(WX5165,WX5142,WX5111);
	and 	XG10392 	(WX5151,WX5142,WX5112);
	and 	XG10393 	(WX3882,WX3849,WX3817);
	and 	XG10394 	(WX3872,WX3849,WX3818);
	and 	XG10395 	(WX3858,WX3849,WX3819);
	and 	XG10396 	(WX2589,WX2556,WX2524);
	and 	XG10397 	(WX2579,WX2556,WX2525);
	and 	XG10398 	(WX2565,WX2556,WX2526);
	and 	XG10399 	(WX1296,WX1263,WX1231);
	and 	XG10400 	(WX1286,WX1263,WX1232);
	and 	XG10401 	(WX1272,WX1263,WX1233);
	nand 	XG10402 	(II2011,II2010,II1986);
	nand 	XG10403 	(II2042,II2041,II2017);
	nand 	XG10404 	(II2073,II2072,II2048);
	nand 	XG10405 	(II2104,II2103,II2079);
	nand 	XG10406 	(II2135,II2134,II2110);
	nand 	XG10407 	(II2166,II2165,II2141);
	nand 	XG10408 	(II2197,II2196,II2172);
	nand 	XG10409 	(II2228,II2227,II2203);
	nand 	XG10410 	(II2259,II2258,II2234);
	nand 	XG10411 	(II2290,II2289,II2265);
	nand 	XG10412 	(II2321,II2320,II2296);
	nand 	XG10413 	(II2352,II2351,II2327);
	nand 	XG10414 	(II2383,II2382,II2358);
	nand 	XG10415 	(II2414,II2413,II2389);
	nand 	XG10416 	(II2445,II2444,II2420);
	nand 	XG10417 	(II2476,II2475,II2451);
	nand 	XG10418 	(II2507,II2506,II2482);
	nand 	XG10419 	(II2538,II2537,II2513);
	nand 	XG10420 	(II2569,II2568,II2544);
	nand 	XG10421 	(II2600,II2599,II2575);
	nand 	XG10422 	(II2631,II2630,II2606);
	nand 	XG10423 	(II2662,II2661,II2637);
	nand 	XG10424 	(II2693,II2692,II2668);
	nand 	XG10425 	(II2724,II2723,II2699);
	nand 	XG10426 	(II2755,II2754,II2730);
	nand 	XG10427 	(II2786,II2785,II2761);
	nand 	XG10428 	(II2817,II2816,II2792);
	nand 	XG10429 	(II2848,II2847,II2823);
	nand 	XG10430 	(II2879,II2878,II2854);
	nand 	XG10431 	(II2910,II2909,II2885);
	nand 	XG10432 	(II2941,II2940,II2916);
	nand 	XG10433 	(II2972,II2971,II2947);
	nand 	XG10434 	(II6016,II6015,II5991);
	nand 	XG10435 	(II6047,II6046,II6022);
	nand 	XG10436 	(II6078,II6077,II6053);
	nand 	XG10437 	(II6109,II6108,II6084);
	nand 	XG10438 	(II6140,II6139,II6115);
	nand 	XG10439 	(II6171,II6170,II6146);
	nand 	XG10440 	(II6202,II6201,II6177);
	nand 	XG10441 	(II6233,II6232,II6208);
	nand 	XG10442 	(II6264,II6263,II6239);
	nand 	XG10443 	(II6295,II6294,II6270);
	nand 	XG10444 	(II6326,II6325,II6301);
	nand 	XG10445 	(II6357,II6356,II6332);
	nand 	XG10446 	(II6388,II6387,II6363);
	nand 	XG10447 	(II6419,II6418,II6394);
	nand 	XG10448 	(II6450,II6449,II6425);
	nand 	XG10449 	(II6481,II6480,II6456);
	nand 	XG10450 	(II6512,II6511,II6487);
	nand 	XG10451 	(II6543,II6542,II6518);
	nand 	XG10452 	(II6574,II6573,II6549);
	nand 	XG10453 	(II6605,II6604,II6580);
	nand 	XG10454 	(II6636,II6635,II6611);
	nand 	XG10455 	(II6667,II6666,II6642);
	nand 	XG10456 	(II6698,II6697,II6673);
	nand 	XG10457 	(II6729,II6728,II6704);
	nand 	XG10458 	(II6760,II6759,II6735);
	nand 	XG10459 	(II6791,II6790,II6766);
	nand 	XG10460 	(II6822,II6821,II6797);
	nand 	XG10461 	(II6853,II6852,II6828);
	nand 	XG10462 	(II6884,II6883,II6859);
	nand 	XG10463 	(II6915,II6914,II6890);
	nand 	XG10464 	(II6946,II6945,II6921);
	nand 	XG10465 	(II6977,II6976,II6952);
	nand 	XG10466 	(II10021,II10020,II9996);
	nand 	XG10467 	(II10052,II10051,II10027);
	nand 	XG10468 	(II10083,II10082,II10058);
	nand 	XG10469 	(II10114,II10113,II10089);
	nand 	XG10470 	(II10145,II10144,II10120);
	nand 	XG10471 	(II10176,II10175,II10151);
	nand 	XG10472 	(II10207,II10206,II10182);
	nand 	XG10473 	(II10238,II10237,II10213);
	nand 	XG10474 	(II10269,II10268,II10244);
	nand 	XG10475 	(II10300,II10299,II10275);
	nand 	XG10476 	(II10331,II10330,II10306);
	nand 	XG10477 	(II10362,II10361,II10337);
	nand 	XG10478 	(II10393,II10392,II10368);
	nand 	XG10479 	(II10424,II10423,II10399);
	nand 	XG10480 	(II10455,II10454,II10430);
	nand 	XG10481 	(II10486,II10485,II10461);
	nand 	XG10482 	(II10517,II10516,II10492);
	nand 	XG10483 	(II10548,II10547,II10523);
	nand 	XG10484 	(II10579,II10578,II10554);
	nand 	XG10485 	(II10610,II10609,II10585);
	nand 	XG10486 	(II10641,II10640,II10616);
	nand 	XG10487 	(II10672,II10671,II10647);
	nand 	XG10488 	(II10703,II10702,II10678);
	nand 	XG10489 	(II10734,II10733,II10709);
	nand 	XG10490 	(II10765,II10764,II10740);
	nand 	XG10491 	(II10796,II10795,II10771);
	nand 	XG10492 	(II10827,II10826,II10802);
	nand 	XG10493 	(II10858,II10857,II10833);
	nand 	XG10494 	(II10889,II10888,II10864);
	nand 	XG10495 	(II10920,II10919,II10895);
	nand 	XG10496 	(II10951,II10950,II10926);
	nand 	XG10497 	(II10982,II10981,II10957);
	nand 	XG10498 	(II14026,II14025,II14001);
	nand 	XG10499 	(II14057,II14056,II14032);
	nand 	XG10500 	(II14088,II14087,II14063);
	nand 	XG10501 	(II14119,II14118,II14094);
	nand 	XG10502 	(II14150,II14149,II14125);
	nand 	XG10503 	(II14181,II14180,II14156);
	nand 	XG10504 	(II14212,II14211,II14187);
	nand 	XG10505 	(II14243,II14242,II14218);
	nand 	XG10506 	(II14274,II14273,II14249);
	nand 	XG10507 	(II14305,II14304,II14280);
	nand 	XG10508 	(II14336,II14335,II14311);
	nand 	XG10509 	(II14367,II14366,II14342);
	nand 	XG10510 	(II14398,II14397,II14373);
	nand 	XG10511 	(II14429,II14428,II14404);
	nand 	XG10512 	(II14460,II14459,II14435);
	nand 	XG10513 	(II14491,II14490,II14466);
	nand 	XG10514 	(II14522,II14521,II14497);
	nand 	XG10515 	(II14553,II14552,II14528);
	nand 	XG10516 	(II14584,II14583,II14559);
	nand 	XG10517 	(II14615,II14614,II14590);
	nand 	XG10518 	(II14646,II14645,II14621);
	nand 	XG10519 	(II14677,II14676,II14652);
	nand 	XG10520 	(II14708,II14707,II14683);
	nand 	XG10521 	(II14739,II14738,II14714);
	nand 	XG10522 	(II14770,II14769,II14745);
	nand 	XG10523 	(II14801,II14800,II14776);
	nand 	XG10524 	(II14832,II14831,II14807);
	nand 	XG10525 	(II14863,II14862,II14838);
	nand 	XG10526 	(II14894,II14893,II14869);
	nand 	XG10527 	(II14925,II14924,II14900);
	nand 	XG10528 	(II14956,II14955,II14931);
	nand 	XG10529 	(II14987,II14986,II14962);
	nand 	XG10530 	(II18031,II18030,II18006);
	nand 	XG10531 	(II18062,II18061,II18037);
	nand 	XG10532 	(II18093,II18092,II18068);
	nand 	XG10533 	(II18124,II18123,II18099);
	nand 	XG10534 	(II18155,II18154,II18130);
	nand 	XG10535 	(II18186,II18185,II18161);
	nand 	XG10536 	(II18217,II18216,II18192);
	nand 	XG10537 	(II18248,II18247,II18223);
	nand 	XG10538 	(II18279,II18278,II18254);
	nand 	XG10539 	(II18310,II18309,II18285);
	nand 	XG10540 	(II18341,II18340,II18316);
	nand 	XG10541 	(II18372,II18371,II18347);
	nand 	XG10542 	(II18403,II18402,II18378);
	nand 	XG10543 	(II18434,II18433,II18409);
	nand 	XG10544 	(II18465,II18464,II18440);
	nand 	XG10545 	(II18496,II18495,II18471);
	nand 	XG10546 	(II18527,II18526,II18502);
	nand 	XG10547 	(II18558,II18557,II18533);
	nand 	XG10548 	(II18589,II18588,II18564);
	nand 	XG10549 	(II18620,II18619,II18595);
	nand 	XG10550 	(II18651,II18650,II18626);
	nand 	XG10551 	(II18682,II18681,II18657);
	nand 	XG10552 	(II18713,II18712,II18688);
	nand 	XG10553 	(II18744,II18743,II18719);
	nand 	XG10554 	(II18775,II18774,II18750);
	nand 	XG10555 	(II18806,II18805,II18781);
	nand 	XG10556 	(II18837,II18836,II18812);
	nand 	XG10557 	(II18868,II18867,II18843);
	nand 	XG10558 	(II18899,II18898,II18874);
	nand 	XG10559 	(II18930,II18929,II18905);
	nand 	XG10560 	(II18961,II18960,II18936);
	nand 	XG10561 	(II18992,II18991,II18967);
	nand 	XG10562 	(II22036,II22035,II22011);
	nand 	XG10563 	(II22067,II22066,II22042);
	nand 	XG10564 	(II22098,II22097,II22073);
	nand 	XG10565 	(II22129,II22128,II22104);
	nand 	XG10566 	(II22160,II22159,II22135);
	nand 	XG10567 	(II22191,II22190,II22166);
	nand 	XG10568 	(II22222,II22221,II22197);
	nand 	XG10569 	(II22253,II22252,II22228);
	nand 	XG10570 	(II22284,II22283,II22259);
	nand 	XG10571 	(II22315,II22314,II22290);
	nand 	XG10572 	(II22346,II22345,II22321);
	nand 	XG10573 	(II22377,II22376,II22352);
	nand 	XG10574 	(II22408,II22407,II22383);
	nand 	XG10575 	(II22439,II22438,II22414);
	nand 	XG10576 	(II22470,II22469,II22445);
	nand 	XG10577 	(II22501,II22500,II22476);
	nand 	XG10578 	(II22532,II22531,II22507);
	nand 	XG10579 	(II22563,II22562,II22538);
	nand 	XG10580 	(II22594,II22593,II22569);
	nand 	XG10581 	(II22625,II22624,II22600);
	nand 	XG10582 	(II22656,II22655,II22631);
	nand 	XG10583 	(II22687,II22686,II22662);
	nand 	XG10584 	(II22718,II22717,II22693);
	nand 	XG10585 	(II22749,II22748,II22724);
	nand 	XG10586 	(II22780,II22779,II22755);
	nand 	XG10587 	(II22811,II22810,II22786);
	nand 	XG10588 	(II22842,II22841,II22817);
	nand 	XG10589 	(II22873,II22872,II22848);
	nand 	XG10590 	(II22904,II22903,II22879);
	nand 	XG10591 	(II22935,II22934,II22910);
	nand 	XG10592 	(II22966,II22965,II22941);
	nand 	XG10593 	(II22997,II22996,II22972);
	nand 	XG10594 	(II26041,II26040,II26016);
	nand 	XG10595 	(II26072,II26071,II26047);
	nand 	XG10596 	(II26103,II26102,II26078);
	nand 	XG10597 	(II26134,II26133,II26109);
	nand 	XG10598 	(II26165,II26164,II26140);
	nand 	XG10599 	(II26196,II26195,II26171);
	nand 	XG10600 	(II26227,II26226,II26202);
	nand 	XG10601 	(II26258,II26257,II26233);
	nand 	XG10602 	(II26289,II26288,II26264);
	nand 	XG10603 	(II26320,II26319,II26295);
	nand 	XG10604 	(II26351,II26350,II26326);
	nand 	XG10605 	(II26382,II26381,II26357);
	nand 	XG10606 	(II26413,II26412,II26388);
	nand 	XG10607 	(II26444,II26443,II26419);
	nand 	XG10608 	(II26475,II26474,II26450);
	nand 	XG10609 	(II26506,II26505,II26481);
	nand 	XG10610 	(II26537,II26536,II26512);
	nand 	XG10611 	(II26568,II26567,II26543);
	nand 	XG10612 	(II26599,II26598,II26574);
	nand 	XG10613 	(II26630,II26629,II26605);
	nand 	XG10614 	(II26661,II26660,II26636);
	nand 	XG10615 	(II26692,II26691,II26667);
	nand 	XG10616 	(II26723,II26722,II26698);
	nand 	XG10617 	(II26754,II26753,II26729);
	nand 	XG10618 	(II26785,II26784,II26760);
	nand 	XG10619 	(II26816,II26815,II26791);
	nand 	XG10620 	(II26847,II26846,II26822);
	nand 	XG10621 	(II26878,II26877,II26853);
	nand 	XG10622 	(II26909,II26908,II26884);
	nand 	XG10623 	(II26940,II26939,II26915);
	nand 	XG10624 	(II26971,II26970,II26946);
	nand 	XG10625 	(II27002,II27001,II26977);
	nand 	XG10626 	(II30046,II30045,II30021);
	nand 	XG10627 	(II30077,II30076,II30052);
	nand 	XG10628 	(II30108,II30107,II30083);
	nand 	XG10629 	(II30139,II30138,II30114);
	nand 	XG10630 	(II30170,II30169,II30145);
	nand 	XG10631 	(II30201,II30200,II30176);
	nand 	XG10632 	(II30232,II30231,II30207);
	nand 	XG10633 	(II30263,II30262,II30238);
	nand 	XG10634 	(II30294,II30293,II30269);
	nand 	XG10635 	(II30325,II30324,II30300);
	nand 	XG10636 	(II30356,II30355,II30331);
	nand 	XG10637 	(II30387,II30386,II30362);
	nand 	XG10638 	(II30418,II30417,II30393);
	nand 	XG10639 	(II30449,II30448,II30424);
	nand 	XG10640 	(II30480,II30479,II30455);
	nand 	XG10641 	(II30511,II30510,II30486);
	nand 	XG10642 	(II30542,II30541,II30517);
	nand 	XG10643 	(II30573,II30572,II30548);
	nand 	XG10644 	(II30604,II30603,II30579);
	nand 	XG10645 	(II30635,II30634,II30610);
	nand 	XG10646 	(II30666,II30665,II30641);
	nand 	XG10647 	(II30697,II30696,II30672);
	nand 	XG10648 	(II30728,II30727,II30703);
	nand 	XG10649 	(II30759,II30758,II30734);
	nand 	XG10650 	(II30790,II30789,II30765);
	nand 	XG10651 	(II30821,II30820,II30796);
	nand 	XG10652 	(II30852,II30851,II30827);
	nand 	XG10653 	(II30883,II30882,II30858);
	nand 	XG10654 	(II30914,II30913,II30889);
	nand 	XG10655 	(II30945,II30944,II30920);
	nand 	XG10656 	(II30976,II30975,II30951);
	nand 	XG10657 	(II31007,II31006,II30982);
	nand 	XG10658 	(II34051,II34050,II34026);
	nand 	XG10659 	(II34082,II34081,II34057);
	nand 	XG10660 	(II34113,II34112,II34088);
	nand 	XG10661 	(II34144,II34143,II34119);
	nand 	XG10662 	(II34175,II34174,II34150);
	nand 	XG10663 	(II34206,II34205,II34181);
	nand 	XG10664 	(II34237,II34236,II34212);
	nand 	XG10665 	(II34268,II34267,II34243);
	nand 	XG10666 	(II34299,II34298,II34274);
	nand 	XG10667 	(II34330,II34329,II34305);
	nand 	XG10668 	(II34361,II34360,II34336);
	nand 	XG10669 	(II34392,II34391,II34367);
	nand 	XG10670 	(II34423,II34422,II34398);
	nand 	XG10671 	(II34454,II34453,II34429);
	nand 	XG10672 	(II34485,II34484,II34460);
	nand 	XG10673 	(II34516,II34515,II34491);
	nand 	XG10674 	(II34547,II34546,II34522);
	nand 	XG10675 	(II34578,II34577,II34553);
	nand 	XG10676 	(II34609,II34608,II34584);
	nand 	XG10677 	(II34640,II34639,II34615);
	nand 	XG10678 	(II34671,II34670,II34646);
	nand 	XG10679 	(II34702,II34701,II34677);
	nand 	XG10680 	(II34733,II34732,II34708);
	nand 	XG10681 	(II34764,II34763,II34739);
	nand 	XG10682 	(II34795,II34794,II34770);
	nand 	XG10683 	(II34826,II34825,II34801);
	nand 	XG10684 	(II34857,II34856,II34832);
	nand 	XG10685 	(II34888,II34887,II34863);
	nand 	XG10686 	(II34919,II34918,II34894);
	nand 	XG10687 	(II34950,II34949,II34925);
	nand 	XG10688 	(II34981,II34980,II34956);
	nand 	XG10689 	(II35012,II35011,II34987);
	nand 	XG10690 	(II35013,II35011,II35003);
	nand 	XG10691 	(II34982,II34980,II34972);
	nand 	XG10692 	(II34951,II34949,II34941);
	nand 	XG10693 	(II34920,II34918,II34910);
	nand 	XG10694 	(II34889,II34887,II34879);
	nand 	XG10695 	(II34858,II34856,II34848);
	nand 	XG10696 	(II34827,II34825,II34817);
	nand 	XG10697 	(II34796,II34794,II34786);
	nand 	XG10698 	(II34765,II34763,II34755);
	nand 	XG10699 	(II34734,II34732,II34724);
	nand 	XG10700 	(II34703,II34701,II34693);
	nand 	XG10701 	(II34672,II34670,II34662);
	nand 	XG10702 	(II34641,II34639,II34631);
	nand 	XG10703 	(II34610,II34608,II34600);
	nand 	XG10704 	(II34579,II34577,II34569);
	nand 	XG10705 	(II34548,II34546,II34538);
	nand 	XG10706 	(II34517,II34515,II34507);
	nand 	XG10707 	(II34486,II34484,II34476);
	nand 	XG10708 	(II34455,II34453,II34445);
	nand 	XG10709 	(II34424,II34422,II34414);
	nand 	XG10710 	(II34393,II34391,II34383);
	nand 	XG10711 	(II34362,II34360,II34352);
	nand 	XG10712 	(II34331,II34329,II34321);
	nand 	XG10713 	(II34300,II34298,II34290);
	nand 	XG10714 	(II34269,II34267,II34259);
	nand 	XG10715 	(II34238,II34236,II34228);
	nand 	XG10716 	(II34207,II34205,II34197);
	nand 	XG10717 	(II34176,II34174,II34166);
	nand 	XG10718 	(II34145,II34143,II34135);
	nand 	XG10719 	(II34114,II34112,II34104);
	nand 	XG10720 	(II34083,II34081,II34073);
	nand 	XG10721 	(II34052,II34050,II34042);
	nand 	XG10722 	(II31008,II31006,II30998);
	nand 	XG10723 	(II30977,II30975,II30967);
	nand 	XG10724 	(II30946,II30944,II30936);
	nand 	XG10725 	(II30915,II30913,II30905);
	nand 	XG10726 	(II30884,II30882,II30874);
	nand 	XG10727 	(II30853,II30851,II30843);
	nand 	XG10728 	(II30822,II30820,II30812);
	nand 	XG10729 	(II30791,II30789,II30781);
	nand 	XG10730 	(II30760,II30758,II30750);
	nand 	XG10731 	(II30729,II30727,II30719);
	nand 	XG10732 	(II30698,II30696,II30688);
	nand 	XG10733 	(II30667,II30665,II30657);
	nand 	XG10734 	(II30636,II30634,II30626);
	nand 	XG10735 	(II30605,II30603,II30595);
	nand 	XG10736 	(II30574,II30572,II30564);
	nand 	XG10737 	(II30543,II30541,II30533);
	nand 	XG10738 	(II30512,II30510,II30502);
	nand 	XG10739 	(II30481,II30479,II30471);
	nand 	XG10740 	(II30450,II30448,II30440);
	nand 	XG10741 	(II30419,II30417,II30409);
	nand 	XG10742 	(II30388,II30386,II30378);
	nand 	XG10743 	(II30357,II30355,II30347);
	nand 	XG10744 	(II30326,II30324,II30316);
	nand 	XG10745 	(II30295,II30293,II30285);
	nand 	XG10746 	(II30264,II30262,II30254);
	nand 	XG10747 	(II30233,II30231,II30223);
	nand 	XG10748 	(II30202,II30200,II30192);
	nand 	XG10749 	(II30171,II30169,II30161);
	nand 	XG10750 	(II30140,II30138,II30130);
	nand 	XG10751 	(II30109,II30107,II30099);
	nand 	XG10752 	(II30078,II30076,II30068);
	nand 	XG10753 	(II30047,II30045,II30037);
	nand 	XG10754 	(II27003,II27001,II26993);
	nand 	XG10755 	(II26972,II26970,II26962);
	nand 	XG10756 	(II26941,II26939,II26931);
	nand 	XG10757 	(II26910,II26908,II26900);
	nand 	XG10758 	(II26879,II26877,II26869);
	nand 	XG10759 	(II26848,II26846,II26838);
	nand 	XG10760 	(II26817,II26815,II26807);
	nand 	XG10761 	(II26786,II26784,II26776);
	nand 	XG10762 	(II26755,II26753,II26745);
	nand 	XG10763 	(II26724,II26722,II26714);
	nand 	XG10764 	(II26693,II26691,II26683);
	nand 	XG10765 	(II26662,II26660,II26652);
	nand 	XG10766 	(II26631,II26629,II26621);
	nand 	XG10767 	(II26600,II26598,II26590);
	nand 	XG10768 	(II26569,II26567,II26559);
	nand 	XG10769 	(II26538,II26536,II26528);
	nand 	XG10770 	(II26507,II26505,II26497);
	nand 	XG10771 	(II26476,II26474,II26466);
	nand 	XG10772 	(II26445,II26443,II26435);
	nand 	XG10773 	(II26414,II26412,II26404);
	nand 	XG10774 	(II26383,II26381,II26373);
	nand 	XG10775 	(II26352,II26350,II26342);
	nand 	XG10776 	(II26321,II26319,II26311);
	nand 	XG10777 	(II26290,II26288,II26280);
	nand 	XG10778 	(II26259,II26257,II26249);
	nand 	XG10779 	(II26228,II26226,II26218);
	nand 	XG10780 	(II26197,II26195,II26187);
	nand 	XG10781 	(II26166,II26164,II26156);
	nand 	XG10782 	(II26135,II26133,II26125);
	nand 	XG10783 	(II26104,II26102,II26094);
	nand 	XG10784 	(II26073,II26071,II26063);
	nand 	XG10785 	(II26042,II26040,II26032);
	nand 	XG10786 	(II22998,II22996,II22988);
	nand 	XG10787 	(II22967,II22965,II22957);
	nand 	XG10788 	(II22936,II22934,II22926);
	nand 	XG10789 	(II22905,II22903,II22895);
	nand 	XG10790 	(II22874,II22872,II22864);
	nand 	XG10791 	(II22843,II22841,II22833);
	nand 	XG10792 	(II22812,II22810,II22802);
	nand 	XG10793 	(II22781,II22779,II22771);
	nand 	XG10794 	(II22750,II22748,II22740);
	nand 	XG10795 	(II22719,II22717,II22709);
	nand 	XG10796 	(II22688,II22686,II22678);
	nand 	XG10797 	(II22657,II22655,II22647);
	nand 	XG10798 	(II22626,II22624,II22616);
	nand 	XG10799 	(II22595,II22593,II22585);
	nand 	XG10800 	(II22564,II22562,II22554);
	nand 	XG10801 	(II22533,II22531,II22523);
	nand 	XG10802 	(II22502,II22500,II22492);
	nand 	XG10803 	(II22471,II22469,II22461);
	nand 	XG10804 	(II22440,II22438,II22430);
	nand 	XG10805 	(II22409,II22407,II22399);
	nand 	XG10806 	(II22378,II22376,II22368);
	nand 	XG10807 	(II22347,II22345,II22337);
	nand 	XG10808 	(II22316,II22314,II22306);
	nand 	XG10809 	(II22285,II22283,II22275);
	nand 	XG10810 	(II22254,II22252,II22244);
	nand 	XG10811 	(II22223,II22221,II22213);
	nand 	XG10812 	(II22192,II22190,II22182);
	nand 	XG10813 	(II22161,II22159,II22151);
	nand 	XG10814 	(II22130,II22128,II22120);
	nand 	XG10815 	(II22099,II22097,II22089);
	nand 	XG10816 	(II22068,II22066,II22058);
	nand 	XG10817 	(II22037,II22035,II22027);
	nand 	XG10818 	(II18993,II18991,II18983);
	nand 	XG10819 	(II18962,II18960,II18952);
	nand 	XG10820 	(II18931,II18929,II18921);
	nand 	XG10821 	(II18900,II18898,II18890);
	nand 	XG10822 	(II18869,II18867,II18859);
	nand 	XG10823 	(II18838,II18836,II18828);
	nand 	XG10824 	(II18807,II18805,II18797);
	nand 	XG10825 	(II18776,II18774,II18766);
	nand 	XG10826 	(II18745,II18743,II18735);
	nand 	XG10827 	(II18714,II18712,II18704);
	nand 	XG10828 	(II18683,II18681,II18673);
	nand 	XG10829 	(II18652,II18650,II18642);
	nand 	XG10830 	(II18621,II18619,II18611);
	nand 	XG10831 	(II18590,II18588,II18580);
	nand 	XG10832 	(II18559,II18557,II18549);
	nand 	XG10833 	(II18528,II18526,II18518);
	nand 	XG10834 	(II18497,II18495,II18487);
	nand 	XG10835 	(II18466,II18464,II18456);
	nand 	XG10836 	(II18435,II18433,II18425);
	nand 	XG10837 	(II18404,II18402,II18394);
	nand 	XG10838 	(II18373,II18371,II18363);
	nand 	XG10839 	(II18342,II18340,II18332);
	nand 	XG10840 	(II18311,II18309,II18301);
	nand 	XG10841 	(II18280,II18278,II18270);
	nand 	XG10842 	(II18249,II18247,II18239);
	nand 	XG10843 	(II18218,II18216,II18208);
	nand 	XG10844 	(II18187,II18185,II18177);
	nand 	XG10845 	(II18156,II18154,II18146);
	nand 	XG10846 	(II18125,II18123,II18115);
	nand 	XG10847 	(II18094,II18092,II18084);
	nand 	XG10848 	(II18063,II18061,II18053);
	nand 	XG10849 	(II18032,II18030,II18022);
	nand 	XG10850 	(II14988,II14986,II14978);
	nand 	XG10851 	(II14957,II14955,II14947);
	nand 	XG10852 	(II14926,II14924,II14916);
	nand 	XG10853 	(II14895,II14893,II14885);
	nand 	XG10854 	(II14864,II14862,II14854);
	nand 	XG10855 	(II14833,II14831,II14823);
	nand 	XG10856 	(II14802,II14800,II14792);
	nand 	XG10857 	(II14771,II14769,II14761);
	nand 	XG10858 	(II14740,II14738,II14730);
	nand 	XG10859 	(II14709,II14707,II14699);
	nand 	XG10860 	(II14678,II14676,II14668);
	nand 	XG10861 	(II14647,II14645,II14637);
	nand 	XG10862 	(II14616,II14614,II14606);
	nand 	XG10863 	(II14585,II14583,II14575);
	nand 	XG10864 	(II14554,II14552,II14544);
	nand 	XG10865 	(II14523,II14521,II14513);
	nand 	XG10866 	(II14492,II14490,II14482);
	nand 	XG10867 	(II14461,II14459,II14451);
	nand 	XG10868 	(II14430,II14428,II14420);
	nand 	XG10869 	(II14399,II14397,II14389);
	nand 	XG10870 	(II14368,II14366,II14358);
	nand 	XG10871 	(II14337,II14335,II14327);
	nand 	XG10872 	(II14306,II14304,II14296);
	nand 	XG10873 	(II14275,II14273,II14265);
	nand 	XG10874 	(II14244,II14242,II14234);
	nand 	XG10875 	(II14213,II14211,II14203);
	nand 	XG10876 	(II14182,II14180,II14172);
	nand 	XG10877 	(II14151,II14149,II14141);
	nand 	XG10878 	(II14120,II14118,II14110);
	nand 	XG10879 	(II14089,II14087,II14079);
	nand 	XG10880 	(II14058,II14056,II14048);
	nand 	XG10881 	(II14027,II14025,II14017);
	nand 	XG10882 	(II10983,II10981,II10973);
	nand 	XG10883 	(II10952,II10950,II10942);
	nand 	XG10884 	(II10921,II10919,II10911);
	nand 	XG10885 	(II10890,II10888,II10880);
	nand 	XG10886 	(II10859,II10857,II10849);
	nand 	XG10887 	(II10828,II10826,II10818);
	nand 	XG10888 	(II10797,II10795,II10787);
	nand 	XG10889 	(II10766,II10764,II10756);
	nand 	XG10890 	(II10735,II10733,II10725);
	nand 	XG10891 	(II10704,II10702,II10694);
	nand 	XG10892 	(II10673,II10671,II10663);
	nand 	XG10893 	(II10642,II10640,II10632);
	nand 	XG10894 	(II10611,II10609,II10601);
	nand 	XG10895 	(II10580,II10578,II10570);
	nand 	XG10896 	(II10549,II10547,II10539);
	nand 	XG10897 	(II10518,II10516,II10508);
	nand 	XG10898 	(II10487,II10485,II10477);
	nand 	XG10899 	(II10456,II10454,II10446);
	nand 	XG10900 	(II10425,II10423,II10415);
	nand 	XG10901 	(II10394,II10392,II10384);
	nand 	XG10902 	(II10363,II10361,II10353);
	nand 	XG10903 	(II10332,II10330,II10322);
	nand 	XG10904 	(II10301,II10299,II10291);
	nand 	XG10905 	(II10270,II10268,II10260);
	nand 	XG10906 	(II10239,II10237,II10229);
	nand 	XG10907 	(II10208,II10206,II10198);
	nand 	XG10908 	(II10177,II10175,II10167);
	nand 	XG10909 	(II10146,II10144,II10136);
	nand 	XG10910 	(II10115,II10113,II10105);
	nand 	XG10911 	(II10084,II10082,II10074);
	nand 	XG10912 	(II10053,II10051,II10043);
	nand 	XG10913 	(II10022,II10020,II10012);
	nand 	XG10914 	(II6978,II6976,II6968);
	nand 	XG10915 	(II6947,II6945,II6937);
	nand 	XG10916 	(II6916,II6914,II6906);
	nand 	XG10917 	(II6885,II6883,II6875);
	nand 	XG10918 	(II6854,II6852,II6844);
	nand 	XG10919 	(II6823,II6821,II6813);
	nand 	XG10920 	(II6792,II6790,II6782);
	nand 	XG10921 	(II6761,II6759,II6751);
	nand 	XG10922 	(II6730,II6728,II6720);
	nand 	XG10923 	(II6699,II6697,II6689);
	nand 	XG10924 	(II6668,II6666,II6658);
	nand 	XG10925 	(II6637,II6635,II6627);
	nand 	XG10926 	(II6606,II6604,II6596);
	nand 	XG10927 	(II6575,II6573,II6565);
	nand 	XG10928 	(II6544,II6542,II6534);
	nand 	XG10929 	(II6513,II6511,II6503);
	nand 	XG10930 	(II6482,II6480,II6472);
	nand 	XG10931 	(II6451,II6449,II6441);
	nand 	XG10932 	(II6420,II6418,II6410);
	nand 	XG10933 	(II6389,II6387,II6379);
	nand 	XG10934 	(II6358,II6356,II6348);
	nand 	XG10935 	(II6327,II6325,II6317);
	nand 	XG10936 	(II6296,II6294,II6286);
	nand 	XG10937 	(II6265,II6263,II6255);
	nand 	XG10938 	(II6234,II6232,II6224);
	nand 	XG10939 	(II6203,II6201,II6193);
	nand 	XG10940 	(II6172,II6170,II6162);
	nand 	XG10941 	(II6141,II6139,II6131);
	nand 	XG10942 	(II6110,II6108,II6100);
	nand 	XG10943 	(II6079,II6077,II6069);
	nand 	XG10944 	(II6048,II6046,II6038);
	nand 	XG10945 	(II6017,II6015,II6007);
	nand 	XG10946 	(II2973,II2971,II2963);
	nand 	XG10947 	(II2942,II2940,II2932);
	nand 	XG10948 	(II2911,II2909,II2901);
	nand 	XG10949 	(II2880,II2878,II2870);
	nand 	XG10950 	(II2849,II2847,II2839);
	nand 	XG10951 	(II2818,II2816,II2808);
	nand 	XG10952 	(II2787,II2785,II2777);
	nand 	XG10953 	(II2756,II2754,II2746);
	nand 	XG10954 	(II2725,II2723,II2715);
	nand 	XG10955 	(II2694,II2692,II2684);
	nand 	XG10956 	(II2663,II2661,II2653);
	nand 	XG10957 	(II2632,II2630,II2622);
	nand 	XG10958 	(II2601,II2599,II2591);
	nand 	XG10959 	(II2570,II2568,II2560);
	nand 	XG10960 	(II2539,II2537,II2529);
	nand 	XG10961 	(II2508,II2506,II2498);
	nand 	XG10962 	(II2477,II2475,II2467);
	nand 	XG10963 	(II2446,II2444,II2436);
	nand 	XG10964 	(II2415,II2413,II2405);
	nand 	XG10965 	(II2384,II2382,II2374);
	nand 	XG10966 	(II2353,II2351,II2343);
	nand 	XG10967 	(II2322,II2320,II2312);
	nand 	XG10968 	(II2291,II2289,II2281);
	nand 	XG10969 	(II2260,II2258,II2250);
	nand 	XG10970 	(II2229,II2227,II2219);
	nand 	XG10971 	(II2198,II2196,II2188);
	nand 	XG10972 	(II2167,II2165,II2157);
	nand 	XG10973 	(II2136,II2134,II2126);
	nand 	XG10974 	(II2105,II2103,II2095);
	nand 	XG10975 	(II2074,II2072,II2064);
	nand 	XG10976 	(II2043,II2041,II2033);
	nand 	XG10977 	(II2012,II2010,II2002);
	nand 	XG10978 	(WX11275,II35013,II35012);
	nand 	XG10979 	(WX11274,II34982,II34981);
	nand 	XG10980 	(WX11273,II34951,II34950);
	nand 	XG10981 	(WX11272,II34920,II34919);
	nand 	XG10982 	(WX11271,II34889,II34888);
	nand 	XG10983 	(WX11270,II34858,II34857);
	nand 	XG10984 	(WX11269,II34827,II34826);
	nand 	XG10985 	(WX11268,II34796,II34795);
	nand 	XG10986 	(WX11267,II34765,II34764);
	nand 	XG10987 	(WX11266,II34734,II34733);
	nand 	XG10988 	(WX11265,II34703,II34702);
	nand 	XG10989 	(WX11264,II34672,II34671);
	nand 	XG10990 	(WX11263,II34641,II34640);
	nand 	XG10991 	(WX11262,II34610,II34609);
	nand 	XG10992 	(WX11261,II34579,II34578);
	nand 	XG10993 	(WX11260,II34548,II34547);
	nand 	XG10994 	(WX11259,II34517,II34516);
	nand 	XG10995 	(WX11258,II34486,II34485);
	nand 	XG10996 	(WX11257,II34455,II34454);
	nand 	XG10997 	(WX11256,II34424,II34423);
	nand 	XG10998 	(WX11255,II34393,II34392);
	nand 	XG10999 	(WX11254,II34362,II34361);
	nand 	XG11000 	(WX11253,II34331,II34330);
	nand 	XG11001 	(WX11252,II34300,II34299);
	nand 	XG11002 	(WX11251,II34269,II34268);
	nand 	XG11003 	(WX11250,II34238,II34237);
	nand 	XG11004 	(WX11249,II34207,II34206);
	nand 	XG11005 	(WX11248,II34176,II34175);
	nand 	XG11006 	(WX11247,II34145,II34144);
	nand 	XG11007 	(WX11246,II34114,II34113);
	nand 	XG11008 	(WX11245,II34083,II34082);
	nand 	XG11009 	(WX11244,II34052,II34051);
	nand 	XG11010 	(WX9982,II31008,II31007);
	nand 	XG11011 	(WX9981,II30977,II30976);
	nand 	XG11012 	(WX9980,II30946,II30945);
	nand 	XG11013 	(WX9979,II30915,II30914);
	nand 	XG11014 	(WX9978,II30884,II30883);
	nand 	XG11015 	(WX9977,II30853,II30852);
	nand 	XG11016 	(WX9976,II30822,II30821);
	nand 	XG11017 	(WX9975,II30791,II30790);
	nand 	XG11018 	(WX9974,II30760,II30759);
	nand 	XG11019 	(WX9973,II30729,II30728);
	nand 	XG11020 	(WX9972,II30698,II30697);
	nand 	XG11021 	(WX9971,II30667,II30666);
	nand 	XG11022 	(WX9970,II30636,II30635);
	nand 	XG11023 	(WX9969,II30605,II30604);
	nand 	XG11024 	(WX9968,II30574,II30573);
	nand 	XG11025 	(WX9967,II30543,II30542);
	nand 	XG11026 	(WX9966,II30512,II30511);
	nand 	XG11027 	(WX9965,II30481,II30480);
	nand 	XG11028 	(WX9964,II30450,II30449);
	nand 	XG11029 	(WX9963,II30419,II30418);
	nand 	XG11030 	(WX9962,II30388,II30387);
	nand 	XG11031 	(WX9961,II30357,II30356);
	nand 	XG11032 	(WX9960,II30326,II30325);
	nand 	XG11033 	(WX9959,II30295,II30294);
	nand 	XG11034 	(WX9958,II30264,II30263);
	nand 	XG11035 	(WX9957,II30233,II30232);
	nand 	XG11036 	(WX9956,II30202,II30201);
	nand 	XG11037 	(WX9955,II30171,II30170);
	nand 	XG11038 	(WX9954,II30140,II30139);
	nand 	XG11039 	(WX9953,II30109,II30108);
	nand 	XG11040 	(WX9952,II30078,II30077);
	nand 	XG11041 	(WX9951,II30047,II30046);
	nand 	XG11042 	(WX8689,II27003,II27002);
	nand 	XG11043 	(WX8688,II26972,II26971);
	nand 	XG11044 	(WX8687,II26941,II26940);
	nand 	XG11045 	(WX8686,II26910,II26909);
	nand 	XG11046 	(WX8685,II26879,II26878);
	nand 	XG11047 	(WX8684,II26848,II26847);
	nand 	XG11048 	(WX8683,II26817,II26816);
	nand 	XG11049 	(WX8682,II26786,II26785);
	nand 	XG11050 	(WX8681,II26755,II26754);
	nand 	XG11051 	(WX8680,II26724,II26723);
	nand 	XG11052 	(WX8679,II26693,II26692);
	nand 	XG11053 	(WX8678,II26662,II26661);
	nand 	XG11054 	(WX8677,II26631,II26630);
	nand 	XG11055 	(WX8676,II26600,II26599);
	nand 	XG11056 	(WX8675,II26569,II26568);
	nand 	XG11057 	(WX8674,II26538,II26537);
	nand 	XG11058 	(WX8673,II26507,II26506);
	nand 	XG11059 	(WX8672,II26476,II26475);
	nand 	XG11060 	(WX8671,II26445,II26444);
	nand 	XG11061 	(WX8670,II26414,II26413);
	nand 	XG11062 	(WX8669,II26383,II26382);
	nand 	XG11063 	(WX8668,II26352,II26351);
	nand 	XG11064 	(WX8667,II26321,II26320);
	nand 	XG11065 	(WX8666,II26290,II26289);
	nand 	XG11066 	(WX8665,II26259,II26258);
	nand 	XG11067 	(WX8664,II26228,II26227);
	nand 	XG11068 	(WX8663,II26197,II26196);
	nand 	XG11069 	(WX8662,II26166,II26165);
	nand 	XG11070 	(WX8661,II26135,II26134);
	nand 	XG11071 	(WX8660,II26104,II26103);
	nand 	XG11072 	(WX8659,II26073,II26072);
	nand 	XG11073 	(WX8658,II26042,II26041);
	nand 	XG11074 	(WX7396,II22998,II22997);
	nand 	XG11075 	(WX7395,II22967,II22966);
	nand 	XG11076 	(WX7394,II22936,II22935);
	nand 	XG11077 	(WX7393,II22905,II22904);
	nand 	XG11078 	(WX7392,II22874,II22873);
	nand 	XG11079 	(WX7391,II22843,II22842);
	nand 	XG11080 	(WX7390,II22812,II22811);
	nand 	XG11081 	(WX7389,II22781,II22780);
	nand 	XG11082 	(WX7388,II22750,II22749);
	nand 	XG11083 	(WX7387,II22719,II22718);
	nand 	XG11084 	(WX7386,II22688,II22687);
	nand 	XG11085 	(WX7385,II22657,II22656);
	nand 	XG11086 	(WX7384,II22626,II22625);
	nand 	XG11087 	(WX7383,II22595,II22594);
	nand 	XG11088 	(WX7382,II22564,II22563);
	nand 	XG11089 	(WX7381,II22533,II22532);
	nand 	XG11090 	(WX7380,II22502,II22501);
	nand 	XG11091 	(WX7379,II22471,II22470);
	nand 	XG11092 	(WX7378,II22440,II22439);
	nand 	XG11093 	(WX7377,II22409,II22408);
	nand 	XG11094 	(WX7376,II22378,II22377);
	nand 	XG11095 	(WX7375,II22347,II22346);
	nand 	XG11096 	(WX7374,II22316,II22315);
	nand 	XG11097 	(WX7373,II22285,II22284);
	nand 	XG11098 	(WX7372,II22254,II22253);
	nand 	XG11099 	(WX7371,II22223,II22222);
	nand 	XG11100 	(WX7370,II22192,II22191);
	nand 	XG11101 	(WX7369,II22161,II22160);
	nand 	XG11102 	(WX7368,II22130,II22129);
	nand 	XG11103 	(WX7367,II22099,II22098);
	nand 	XG11104 	(WX7366,II22068,II22067);
	nand 	XG11105 	(WX7365,II22037,II22036);
	nand 	XG11106 	(WX6103,II18993,II18992);
	nand 	XG11107 	(WX6102,II18962,II18961);
	nand 	XG11108 	(WX6101,II18931,II18930);
	nand 	XG11109 	(WX6100,II18900,II18899);
	nand 	XG11110 	(WX6099,II18869,II18868);
	nand 	XG11111 	(WX6098,II18838,II18837);
	nand 	XG11112 	(WX6097,II18807,II18806);
	nand 	XG11113 	(WX6096,II18776,II18775);
	nand 	XG11114 	(WX6095,II18745,II18744);
	nand 	XG11115 	(WX6094,II18714,II18713);
	nand 	XG11116 	(WX6093,II18683,II18682);
	nand 	XG11117 	(WX6092,II18652,II18651);
	nand 	XG11118 	(WX6091,II18621,II18620);
	nand 	XG11119 	(WX6090,II18590,II18589);
	nand 	XG11120 	(WX6089,II18559,II18558);
	nand 	XG11121 	(WX6088,II18528,II18527);
	nand 	XG11122 	(WX6087,II18497,II18496);
	nand 	XG11123 	(WX6086,II18466,II18465);
	nand 	XG11124 	(WX6085,II18435,II18434);
	nand 	XG11125 	(WX6084,II18404,II18403);
	nand 	XG11126 	(WX6083,II18373,II18372);
	nand 	XG11127 	(WX6082,II18342,II18341);
	nand 	XG11128 	(WX6081,II18311,II18310);
	nand 	XG11129 	(WX6080,II18280,II18279);
	nand 	XG11130 	(WX6079,II18249,II18248);
	nand 	XG11131 	(WX6078,II18218,II18217);
	nand 	XG11132 	(WX6077,II18187,II18186);
	nand 	XG11133 	(WX6076,II18156,II18155);
	nand 	XG11134 	(WX6075,II18125,II18124);
	nand 	XG11135 	(WX6074,II18094,II18093);
	nand 	XG11136 	(WX6073,II18063,II18062);
	nand 	XG11137 	(WX6072,II18032,II18031);
	nand 	XG11138 	(WX4810,II14988,II14987);
	nand 	XG11139 	(WX4809,II14957,II14956);
	nand 	XG11140 	(WX4808,II14926,II14925);
	nand 	XG11141 	(WX4807,II14895,II14894);
	nand 	XG11142 	(WX4806,II14864,II14863);
	nand 	XG11143 	(WX4805,II14833,II14832);
	nand 	XG11144 	(WX4804,II14802,II14801);
	nand 	XG11145 	(WX4803,II14771,II14770);
	nand 	XG11146 	(WX4802,II14740,II14739);
	nand 	XG11147 	(WX4801,II14709,II14708);
	nand 	XG11148 	(WX4800,II14678,II14677);
	nand 	XG11149 	(WX4799,II14647,II14646);
	nand 	XG11150 	(WX4798,II14616,II14615);
	nand 	XG11151 	(WX4797,II14585,II14584);
	nand 	XG11152 	(WX4796,II14554,II14553);
	nand 	XG11153 	(WX4795,II14523,II14522);
	nand 	XG11154 	(WX4794,II14492,II14491);
	nand 	XG11155 	(WX4793,II14461,II14460);
	nand 	XG11156 	(WX4792,II14430,II14429);
	nand 	XG11157 	(WX4791,II14399,II14398);
	nand 	XG11158 	(WX4790,II14368,II14367);
	nand 	XG11159 	(WX4789,II14337,II14336);
	nand 	XG11160 	(WX4788,II14306,II14305);
	nand 	XG11161 	(WX4787,II14275,II14274);
	nand 	XG11162 	(WX4786,II14244,II14243);
	nand 	XG11163 	(WX4785,II14213,II14212);
	nand 	XG11164 	(WX4784,II14182,II14181);
	nand 	XG11165 	(WX4783,II14151,II14150);
	nand 	XG11166 	(WX4782,II14120,II14119);
	nand 	XG11167 	(WX4781,II14089,II14088);
	nand 	XG11168 	(WX4780,II14058,II14057);
	nand 	XG11169 	(WX4779,II14027,II14026);
	nand 	XG11170 	(WX3517,II10983,II10982);
	nand 	XG11171 	(WX3516,II10952,II10951);
	nand 	XG11172 	(WX3515,II10921,II10920);
	nand 	XG11173 	(WX3514,II10890,II10889);
	nand 	XG11174 	(WX3513,II10859,II10858);
	nand 	XG11175 	(WX3512,II10828,II10827);
	nand 	XG11176 	(WX3511,II10797,II10796);
	nand 	XG11177 	(WX3510,II10766,II10765);
	nand 	XG11178 	(WX3509,II10735,II10734);
	nand 	XG11179 	(WX3508,II10704,II10703);
	nand 	XG11180 	(WX3507,II10673,II10672);
	nand 	XG11181 	(WX3506,II10642,II10641);
	nand 	XG11182 	(WX3505,II10611,II10610);
	nand 	XG11183 	(WX3504,II10580,II10579);
	nand 	XG11184 	(WX3503,II10549,II10548);
	nand 	XG11185 	(WX3502,II10518,II10517);
	nand 	XG11186 	(WX3501,II10487,II10486);
	nand 	XG11187 	(WX3500,II10456,II10455);
	nand 	XG11188 	(WX3499,II10425,II10424);
	nand 	XG11189 	(WX3498,II10394,II10393);
	nand 	XG11190 	(WX3497,II10363,II10362);
	nand 	XG11191 	(WX3496,II10332,II10331);
	nand 	XG11192 	(WX3495,II10301,II10300);
	nand 	XG11193 	(WX3494,II10270,II10269);
	nand 	XG11194 	(WX3493,II10239,II10238);
	nand 	XG11195 	(WX3492,II10208,II10207);
	nand 	XG11196 	(WX3491,II10177,II10176);
	nand 	XG11197 	(WX3490,II10146,II10145);
	nand 	XG11198 	(WX3489,II10115,II10114);
	nand 	XG11199 	(WX3488,II10084,II10083);
	nand 	XG11200 	(WX3487,II10053,II10052);
	nand 	XG11201 	(WX3486,II10022,II10021);
	nand 	XG11202 	(WX2224,II6978,II6977);
	nand 	XG11203 	(WX2223,II6947,II6946);
	nand 	XG11204 	(WX2222,II6916,II6915);
	nand 	XG11205 	(WX2221,II6885,II6884);
	nand 	XG11206 	(WX2220,II6854,II6853);
	nand 	XG11207 	(WX2219,II6823,II6822);
	nand 	XG11208 	(WX2218,II6792,II6791);
	nand 	XG11209 	(WX2217,II6761,II6760);
	nand 	XG11210 	(WX2216,II6730,II6729);
	nand 	XG11211 	(WX2215,II6699,II6698);
	nand 	XG11212 	(WX2214,II6668,II6667);
	nand 	XG11213 	(WX2213,II6637,II6636);
	nand 	XG11214 	(WX2212,II6606,II6605);
	nand 	XG11215 	(WX2211,II6575,II6574);
	nand 	XG11216 	(WX2210,II6544,II6543);
	nand 	XG11217 	(WX2209,II6513,II6512);
	nand 	XG11218 	(WX2208,II6482,II6481);
	nand 	XG11219 	(WX2207,II6451,II6450);
	nand 	XG11220 	(WX2206,II6420,II6419);
	nand 	XG11221 	(WX2205,II6389,II6388);
	nand 	XG11222 	(WX2204,II6358,II6357);
	nand 	XG11223 	(WX2203,II6327,II6326);
	nand 	XG11224 	(WX2202,II6296,II6295);
	nand 	XG11225 	(WX2201,II6265,II6264);
	nand 	XG11226 	(WX2200,II6234,II6233);
	nand 	XG11227 	(WX2199,II6203,II6202);
	nand 	XG11228 	(WX2198,II6172,II6171);
	nand 	XG11229 	(WX2197,II6141,II6140);
	nand 	XG11230 	(WX2196,II6110,II6109);
	nand 	XG11231 	(WX2195,II6079,II6078);
	nand 	XG11232 	(WX2194,II6048,II6047);
	nand 	XG11233 	(WX2193,II6017,II6016);
	nand 	XG11234 	(WX931,II2973,II2972);
	nand 	XG11235 	(WX930,II2942,II2941);
	nand 	XG11236 	(WX929,II2911,II2910);
	nand 	XG11237 	(WX928,II2880,II2879);
	nand 	XG11238 	(WX927,II2849,II2848);
	nand 	XG11239 	(WX926,II2818,II2817);
	nand 	XG11240 	(WX925,II2787,II2786);
	nand 	XG11241 	(WX924,II2756,II2755);
	nand 	XG11242 	(WX923,II2725,II2724);
	nand 	XG11243 	(WX922,II2694,II2693);
	nand 	XG11244 	(WX921,II2663,II2662);
	nand 	XG11245 	(WX920,II2632,II2631);
	nand 	XG11246 	(WX919,II2601,II2600);
	nand 	XG11247 	(WX918,II2570,II2569);
	nand 	XG11248 	(WX917,II2539,II2538);
	nand 	XG11249 	(WX916,II2508,II2507);
	nand 	XG11250 	(WX915,II2477,II2476);
	nand 	XG11251 	(WX914,II2446,II2445);
	nand 	XG11252 	(WX913,II2415,II2414);
	nand 	XG11253 	(WX912,II2384,II2383);
	nand 	XG11254 	(WX911,II2353,II2352);
	nand 	XG11255 	(WX910,II2322,II2321);
	nand 	XG11256 	(WX909,II2291,II2290);
	nand 	XG11257 	(WX908,II2260,II2259);
	nand 	XG11258 	(WX907,II2229,II2228);
	nand 	XG11259 	(WX906,II2198,II2197);
	nand 	XG11260 	(WX905,II2167,II2166);
	nand 	XG11261 	(WX904,II2136,II2135);
	nand 	XG11262 	(WX903,II2105,II2104);
	nand 	XG11263 	(WX902,II2074,II2073);
	nand 	XG11264 	(WX901,II2043,II2042);
	nand 	XG11265 	(WX900,II2012,II2011);
	not 	XG11266 	(WX964,WX900);
	not 	XG11267 	(WX966,WX901);
	not 	XG11268 	(WX968,WX902);
	not 	XG11269 	(WX970,WX903);
	not 	XG11270 	(WX972,WX904);
	not 	XG11271 	(WX974,WX905);
	not 	XG11272 	(WX976,WX906);
	not 	XG11273 	(WX978,WX907);
	not 	XG11274 	(WX980,WX908);
	not 	XG11275 	(WX982,WX909);
	not 	XG11276 	(WX984,WX910);
	not 	XG11277 	(WX986,WX911);
	not 	XG11278 	(WX988,WX912);
	not 	XG11279 	(WX990,WX913);
	not 	XG11280 	(WX992,WX914);
	not 	XG11281 	(WX994,WX915);
	not 	XG11282 	(WX932,WX916);
	not 	XG11283 	(WX934,WX917);
	not 	XG11284 	(WX936,WX918);
	not 	XG11285 	(WX938,WX919);
	not 	XG11286 	(WX940,WX920);
	not 	XG11287 	(WX942,WX921);
	not 	XG11288 	(WX944,WX922);
	not 	XG11289 	(WX946,WX923);
	not 	XG11290 	(WX948,WX924);
	not 	XG11291 	(WX950,WX925);
	not 	XG11292 	(WX952,WX926);
	not 	XG11293 	(WX954,WX927);
	not 	XG11294 	(WX956,WX928);
	not 	XG11295 	(WX958,WX929);
	not 	XG11296 	(WX960,WX930);
	not 	XG11297 	(WX962,WX931);
	not 	XG11298 	(WX2257,WX2193);
	not 	XG11299 	(WX2259,WX2194);
	not 	XG11300 	(WX2261,WX2195);
	not 	XG11301 	(WX2263,WX2196);
	not 	XG11302 	(WX2265,WX2197);
	not 	XG11303 	(WX2267,WX2198);
	not 	XG11304 	(WX2269,WX2199);
	not 	XG11305 	(WX2271,WX2200);
	not 	XG11306 	(WX2273,WX2201);
	not 	XG11307 	(WX2275,WX2202);
	not 	XG11308 	(WX2277,WX2203);
	not 	XG11309 	(WX2279,WX2204);
	not 	XG11310 	(WX2281,WX2205);
	not 	XG11311 	(WX2283,WX2206);
	not 	XG11312 	(WX2285,WX2207);
	not 	XG11313 	(WX2287,WX2208);
	not 	XG11314 	(WX2225,WX2209);
	not 	XG11315 	(WX2227,WX2210);
	not 	XG11316 	(WX2229,WX2211);
	not 	XG11317 	(WX2231,WX2212);
	not 	XG11318 	(WX2233,WX2213);
	not 	XG11319 	(WX2235,WX2214);
	not 	XG11320 	(WX2237,WX2215);
	not 	XG11321 	(WX2239,WX2216);
	not 	XG11322 	(WX2241,WX2217);
	not 	XG11323 	(WX2243,WX2218);
	not 	XG11324 	(WX2245,WX2219);
	not 	XG11325 	(WX2247,WX2220);
	not 	XG11326 	(WX2249,WX2221);
	not 	XG11327 	(WX2251,WX2222);
	not 	XG11328 	(WX2253,WX2223);
	not 	XG11329 	(WX2255,WX2224);
	not 	XG11330 	(WX3550,WX3486);
	not 	XG11331 	(WX3552,WX3487);
	not 	XG11332 	(WX3554,WX3488);
	not 	XG11333 	(WX3556,WX3489);
	not 	XG11334 	(WX3558,WX3490);
	not 	XG11335 	(WX3560,WX3491);
	not 	XG11336 	(WX3562,WX3492);
	not 	XG11337 	(WX3564,WX3493);
	not 	XG11338 	(WX3566,WX3494);
	not 	XG11339 	(WX3568,WX3495);
	not 	XG11340 	(WX3570,WX3496);
	not 	XG11341 	(WX3572,WX3497);
	not 	XG11342 	(WX3574,WX3498);
	not 	XG11343 	(WX3576,WX3499);
	not 	XG11344 	(WX3578,WX3500);
	not 	XG11345 	(WX3580,WX3501);
	not 	XG11346 	(WX3518,WX3502);
	not 	XG11347 	(WX3520,WX3503);
	not 	XG11348 	(WX3522,WX3504);
	not 	XG11349 	(WX3524,WX3505);
	not 	XG11350 	(WX3526,WX3506);
	not 	XG11351 	(WX3528,WX3507);
	not 	XG11352 	(WX3530,WX3508);
	not 	XG11353 	(WX3532,WX3509);
	not 	XG11354 	(WX3534,WX3510);
	not 	XG11355 	(WX3536,WX3511);
	not 	XG11356 	(WX3538,WX3512);
	not 	XG11357 	(WX3540,WX3513);
	not 	XG11358 	(WX3542,WX3514);
	not 	XG11359 	(WX3544,WX3515);
	not 	XG11360 	(WX3546,WX3516);
	not 	XG11361 	(WX3548,WX3517);
	not 	XG11362 	(WX4843,WX4779);
	not 	XG11363 	(WX4845,WX4780);
	not 	XG11364 	(WX4847,WX4781);
	not 	XG11365 	(WX4849,WX4782);
	not 	XG11366 	(WX4851,WX4783);
	not 	XG11367 	(WX4853,WX4784);
	not 	XG11368 	(WX4855,WX4785);
	not 	XG11369 	(WX4857,WX4786);
	not 	XG11370 	(WX4859,WX4787);
	not 	XG11371 	(WX4861,WX4788);
	not 	XG11372 	(WX4863,WX4789);
	not 	XG11373 	(WX4865,WX4790);
	not 	XG11374 	(WX4867,WX4791);
	not 	XG11375 	(WX4869,WX4792);
	not 	XG11376 	(WX4871,WX4793);
	not 	XG11377 	(WX4873,WX4794);
	not 	XG11378 	(WX4811,WX4795);
	not 	XG11379 	(WX4813,WX4796);
	not 	XG11380 	(WX4815,WX4797);
	not 	XG11381 	(WX4817,WX4798);
	not 	XG11382 	(WX4819,WX4799);
	not 	XG11383 	(WX4821,WX4800);
	not 	XG11384 	(WX4823,WX4801);
	not 	XG11385 	(WX4825,WX4802);
	not 	XG11386 	(WX4827,WX4803);
	not 	XG11387 	(WX4829,WX4804);
	not 	XG11388 	(WX4831,WX4805);
	not 	XG11389 	(WX4833,WX4806);
	not 	XG11390 	(WX4835,WX4807);
	not 	XG11391 	(WX4837,WX4808);
	not 	XG11392 	(WX4839,WX4809);
	not 	XG11393 	(WX4841,WX4810);
	not 	XG11394 	(WX6136,WX6072);
	not 	XG11395 	(WX6138,WX6073);
	not 	XG11396 	(WX6140,WX6074);
	not 	XG11397 	(WX6142,WX6075);
	not 	XG11398 	(WX6144,WX6076);
	not 	XG11399 	(WX6146,WX6077);
	not 	XG11400 	(WX6148,WX6078);
	not 	XG11401 	(WX6150,WX6079);
	not 	XG11402 	(WX6152,WX6080);
	not 	XG11403 	(WX6154,WX6081);
	not 	XG11404 	(WX6156,WX6082);
	not 	XG11405 	(WX6158,WX6083);
	not 	XG11406 	(WX6160,WX6084);
	not 	XG11407 	(WX6162,WX6085);
	not 	XG11408 	(WX6164,WX6086);
	not 	XG11409 	(WX6166,WX6087);
	not 	XG11410 	(WX6104,WX6088);
	not 	XG11411 	(WX6106,WX6089);
	not 	XG11412 	(WX6108,WX6090);
	not 	XG11413 	(WX6110,WX6091);
	not 	XG11414 	(WX6112,WX6092);
	not 	XG11415 	(WX6114,WX6093);
	not 	XG11416 	(WX6116,WX6094);
	not 	XG11417 	(WX6118,WX6095);
	not 	XG11418 	(WX6120,WX6096);
	not 	XG11419 	(WX6122,WX6097);
	not 	XG11420 	(WX6124,WX6098);
	not 	XG11421 	(WX6126,WX6099);
	not 	XG11422 	(WX6128,WX6100);
	not 	XG11423 	(WX6130,WX6101);
	not 	XG11424 	(WX6132,WX6102);
	not 	XG11425 	(WX6134,WX6103);
	not 	XG11426 	(WX7429,WX7365);
	not 	XG11427 	(WX7431,WX7366);
	not 	XG11428 	(WX7433,WX7367);
	not 	XG11429 	(WX7435,WX7368);
	not 	XG11430 	(WX7437,WX7369);
	not 	XG11431 	(WX7439,WX7370);
	not 	XG11432 	(WX7441,WX7371);
	not 	XG11433 	(WX7443,WX7372);
	not 	XG11434 	(WX7445,WX7373);
	not 	XG11435 	(WX7447,WX7374);
	not 	XG11436 	(WX7449,WX7375);
	not 	XG11437 	(WX7451,WX7376);
	not 	XG11438 	(WX7453,WX7377);
	not 	XG11439 	(WX7455,WX7378);
	not 	XG11440 	(WX7457,WX7379);
	not 	XG11441 	(WX7459,WX7380);
	not 	XG11442 	(WX7397,WX7381);
	not 	XG11443 	(WX7399,WX7382);
	not 	XG11444 	(WX7401,WX7383);
	not 	XG11445 	(WX7403,WX7384);
	not 	XG11446 	(WX7405,WX7385);
	not 	XG11447 	(WX7407,WX7386);
	not 	XG11448 	(WX7409,WX7387);
	not 	XG11449 	(WX7411,WX7388);
	not 	XG11450 	(WX7413,WX7389);
	not 	XG11451 	(WX7415,WX7390);
	not 	XG11452 	(WX7417,WX7391);
	not 	XG11453 	(WX7419,WX7392);
	not 	XG11454 	(WX7421,WX7393);
	not 	XG11455 	(WX7423,WX7394);
	not 	XG11456 	(WX7425,WX7395);
	not 	XG11457 	(WX7427,WX7396);
	not 	XG11458 	(WX8722,WX8658);
	not 	XG11459 	(WX8724,WX8659);
	not 	XG11460 	(WX8726,WX8660);
	not 	XG11461 	(WX8728,WX8661);
	not 	XG11462 	(WX8730,WX8662);
	not 	XG11463 	(WX8732,WX8663);
	not 	XG11464 	(WX8734,WX8664);
	not 	XG11465 	(WX8736,WX8665);
	not 	XG11466 	(WX8738,WX8666);
	not 	XG11467 	(WX8740,WX8667);
	not 	XG11468 	(WX8742,WX8668);
	not 	XG11469 	(WX8744,WX8669);
	not 	XG11470 	(WX8746,WX8670);
	not 	XG11471 	(WX8748,WX8671);
	not 	XG11472 	(WX8750,WX8672);
	not 	XG11473 	(WX8752,WX8673);
	not 	XG11474 	(WX8690,WX8674);
	not 	XG11475 	(WX8692,WX8675);
	not 	XG11476 	(WX8694,WX8676);
	not 	XG11477 	(WX8696,WX8677);
	not 	XG11478 	(WX8698,WX8678);
	not 	XG11479 	(WX8700,WX8679);
	not 	XG11480 	(WX8702,WX8680);
	not 	XG11481 	(WX8704,WX8681);
	not 	XG11482 	(WX8706,WX8682);
	not 	XG11483 	(WX8708,WX8683);
	not 	XG11484 	(WX8710,WX8684);
	not 	XG11485 	(WX8712,WX8685);
	not 	XG11486 	(WX8714,WX8686);
	not 	XG11487 	(WX8716,WX8687);
	not 	XG11488 	(WX8718,WX8688);
	not 	XG11489 	(WX8720,WX8689);
	not 	XG11490 	(WX10015,WX9951);
	not 	XG11491 	(WX10017,WX9952);
	not 	XG11492 	(WX10019,WX9953);
	not 	XG11493 	(WX10021,WX9954);
	not 	XG11494 	(WX10023,WX9955);
	not 	XG11495 	(WX10025,WX9956);
	not 	XG11496 	(WX10027,WX9957);
	not 	XG11497 	(WX10029,WX9958);
	not 	XG11498 	(WX10031,WX9959);
	not 	XG11499 	(WX10033,WX9960);
	not 	XG11500 	(WX10035,WX9961);
	not 	XG11501 	(WX10037,WX9962);
	not 	XG11502 	(WX10039,WX9963);
	not 	XG11503 	(WX10041,WX9964);
	not 	XG11504 	(WX10043,WX9965);
	not 	XG11505 	(WX10045,WX9966);
	not 	XG11506 	(WX9983,WX9967);
	not 	XG11507 	(WX9985,WX9968);
	not 	XG11508 	(WX9987,WX9969);
	not 	XG11509 	(WX9989,WX9970);
	not 	XG11510 	(WX9991,WX9971);
	not 	XG11511 	(WX9993,WX9972);
	not 	XG11512 	(WX9995,WX9973);
	not 	XG11513 	(WX9997,WX9974);
	not 	XG11514 	(WX9999,WX9975);
	not 	XG11515 	(WX10001,WX9976);
	not 	XG11516 	(WX10003,WX9977);
	not 	XG11517 	(WX10005,WX9978);
	not 	XG11518 	(WX10007,WX9979);
	not 	XG11519 	(WX10009,WX9980);
	not 	XG11520 	(WX10011,WX9981);
	not 	XG11521 	(WX10013,WX9982);
	not 	XG11522 	(WX11308,WX11244);
	not 	XG11523 	(WX11310,WX11245);
	not 	XG11524 	(WX11312,WX11246);
	not 	XG11525 	(WX11314,WX11247);
	not 	XG11526 	(WX11316,WX11248);
	not 	XG11527 	(WX11318,WX11249);
	not 	XG11528 	(WX11320,WX11250);
	not 	XG11529 	(WX11322,WX11251);
	not 	XG11530 	(WX11324,WX11252);
	not 	XG11531 	(WX11326,WX11253);
	not 	XG11532 	(WX11328,WX11254);
	not 	XG11533 	(WX11330,WX11255);
	not 	XG11534 	(WX11332,WX11256);
	not 	XG11535 	(WX11334,WX11257);
	not 	XG11536 	(WX11336,WX11258);
	not 	XG11537 	(WX11338,WX11259);
	not 	XG11538 	(WX11276,WX11260);
	not 	XG11539 	(WX11278,WX11261);
	not 	XG11540 	(WX11280,WX11262);
	not 	XG11541 	(WX11282,WX11263);
	not 	XG11542 	(WX11284,WX11264);
	not 	XG11543 	(WX11286,WX11265);
	not 	XG11544 	(WX11288,WX11266);
	not 	XG11545 	(WX11290,WX11267);
	not 	XG11546 	(WX11292,WX11268);
	not 	XG11547 	(WX11294,WX11269);
	not 	XG11548 	(WX11296,WX11270);
	not 	XG11549 	(WX11298,WX11271);
	not 	XG11550 	(WX11300,WX11272);
	not 	XG11551 	(WX11302,WX11273);
	not 	XG11552 	(WX11304,WX11274);
	not 	XG11553 	(WX11306,WX11275);
	not 	XG11554 	(WX11307,WX11306);
	not 	XG11555 	(WX11305,WX11304);
	not 	XG11556 	(WX11303,WX11302);
	not 	XG11557 	(WX11301,WX11300);
	not 	XG11558 	(WX11299,WX11298);
	not 	XG11559 	(WX11297,WX11296);
	not 	XG11560 	(WX11295,WX11294);
	not 	XG11561 	(WX11293,WX11292);
	not 	XG11562 	(WX11291,WX11290);
	not 	XG11563 	(WX11289,WX11288);
	not 	XG11564 	(WX11287,WX11286);
	not 	XG11565 	(WX11285,WX11284);
	not 	XG11566 	(WX11283,WX11282);
	not 	XG11567 	(WX11281,WX11280);
	not 	XG11568 	(WX11279,WX11278);
	not 	XG11569 	(WX11277,WX11276);
	not 	XG11570 	(WX11339,WX11338);
	not 	XG11571 	(WX11337,WX11336);
	not 	XG11572 	(WX11335,WX11334);
	not 	XG11573 	(WX11333,WX11332);
	not 	XG11574 	(WX11331,WX11330);
	not 	XG11575 	(WX11329,WX11328);
	not 	XG11576 	(WX11327,WX11326);
	not 	XG11577 	(WX11325,WX11324);
	not 	XG11578 	(WX11323,WX11322);
	not 	XG11579 	(WX11321,WX11320);
	not 	XG11580 	(WX11319,WX11318);
	not 	XG11581 	(WX11317,WX11316);
	not 	XG11582 	(WX11315,WX11314);
	not 	XG11583 	(WX11313,WX11312);
	not 	XG11584 	(WX11311,WX11310);
	not 	XG11585 	(WX11309,WX11308);
	not 	XG11586 	(WX10014,WX10013);
	not 	XG11587 	(WX10012,WX10011);
	not 	XG11588 	(WX10010,WX10009);
	not 	XG11589 	(WX10008,WX10007);
	not 	XG11590 	(WX10006,WX10005);
	not 	XG11591 	(WX10004,WX10003);
	not 	XG11592 	(WX10002,WX10001);
	not 	XG11593 	(WX10000,WX9999);
	not 	XG11594 	(WX9998,WX9997);
	not 	XG11595 	(WX9996,WX9995);
	not 	XG11596 	(WX9994,WX9993);
	not 	XG11597 	(WX9992,WX9991);
	not 	XG11598 	(WX9990,WX9989);
	not 	XG11599 	(WX9988,WX9987);
	not 	XG11600 	(WX9986,WX9985);
	not 	XG11601 	(WX9984,WX9983);
	not 	XG11602 	(WX10046,WX10045);
	not 	XG11603 	(WX10044,WX10043);
	not 	XG11604 	(WX10042,WX10041);
	not 	XG11605 	(WX10040,WX10039);
	not 	XG11606 	(WX10038,WX10037);
	not 	XG11607 	(WX10036,WX10035);
	not 	XG11608 	(WX10034,WX10033);
	not 	XG11609 	(WX10032,WX10031);
	not 	XG11610 	(WX10030,WX10029);
	not 	XG11611 	(WX10028,WX10027);
	not 	XG11612 	(WX10026,WX10025);
	not 	XG11613 	(WX10024,WX10023);
	not 	XG11614 	(WX10022,WX10021);
	not 	XG11615 	(WX10020,WX10019);
	not 	XG11616 	(WX10018,WX10017);
	not 	XG11617 	(WX10016,WX10015);
	not 	XG11618 	(WX8721,WX8720);
	not 	XG11619 	(WX8719,WX8718);
	not 	XG11620 	(WX8717,WX8716);
	not 	XG11621 	(WX8715,WX8714);
	not 	XG11622 	(WX8713,WX8712);
	not 	XG11623 	(WX8711,WX8710);
	not 	XG11624 	(WX8709,WX8708);
	not 	XG11625 	(WX8707,WX8706);
	not 	XG11626 	(WX8705,WX8704);
	not 	XG11627 	(WX8703,WX8702);
	not 	XG11628 	(WX8701,WX8700);
	not 	XG11629 	(WX8699,WX8698);
	not 	XG11630 	(WX8697,WX8696);
	not 	XG11631 	(WX8695,WX8694);
	not 	XG11632 	(WX8693,WX8692);
	not 	XG11633 	(WX8691,WX8690);
	not 	XG11634 	(WX8753,WX8752);
	not 	XG11635 	(WX8751,WX8750);
	not 	XG11636 	(WX8749,WX8748);
	not 	XG11637 	(WX8747,WX8746);
	not 	XG11638 	(WX8745,WX8744);
	not 	XG11639 	(WX8743,WX8742);
	not 	XG11640 	(WX8741,WX8740);
	not 	XG11641 	(WX8739,WX8738);
	not 	XG11642 	(WX8737,WX8736);
	not 	XG11643 	(WX8735,WX8734);
	not 	XG11644 	(WX8733,WX8732);
	not 	XG11645 	(WX8731,WX8730);
	not 	XG11646 	(WX8729,WX8728);
	not 	XG11647 	(WX8727,WX8726);
	not 	XG11648 	(WX8725,WX8724);
	not 	XG11649 	(WX8723,WX8722);
	not 	XG11650 	(WX7428,WX7427);
	not 	XG11651 	(WX7426,WX7425);
	not 	XG11652 	(WX7424,WX7423);
	not 	XG11653 	(WX7422,WX7421);
	not 	XG11654 	(WX7420,WX7419);
	not 	XG11655 	(WX7418,WX7417);
	not 	XG11656 	(WX7416,WX7415);
	not 	XG11657 	(WX7414,WX7413);
	not 	XG11658 	(WX7412,WX7411);
	not 	XG11659 	(WX7410,WX7409);
	not 	XG11660 	(WX7408,WX7407);
	not 	XG11661 	(WX7406,WX7405);
	not 	XG11662 	(WX7404,WX7403);
	not 	XG11663 	(WX7402,WX7401);
	not 	XG11664 	(WX7400,WX7399);
	not 	XG11665 	(WX7398,WX7397);
	not 	XG11666 	(WX7460,WX7459);
	not 	XG11667 	(WX7458,WX7457);
	not 	XG11668 	(WX7456,WX7455);
	not 	XG11669 	(WX7454,WX7453);
	not 	XG11670 	(WX7452,WX7451);
	not 	XG11671 	(WX7450,WX7449);
	not 	XG11672 	(WX7448,WX7447);
	not 	XG11673 	(WX7446,WX7445);
	not 	XG11674 	(WX7444,WX7443);
	not 	XG11675 	(WX7442,WX7441);
	not 	XG11676 	(WX7440,WX7439);
	not 	XG11677 	(WX7438,WX7437);
	not 	XG11678 	(WX7436,WX7435);
	not 	XG11679 	(WX7434,WX7433);
	not 	XG11680 	(WX7432,WX7431);
	not 	XG11681 	(WX7430,WX7429);
	not 	XG11682 	(WX6135,WX6134);
	not 	XG11683 	(WX6133,WX6132);
	not 	XG11684 	(WX6131,WX6130);
	not 	XG11685 	(WX6129,WX6128);
	not 	XG11686 	(WX6127,WX6126);
	not 	XG11687 	(WX6125,WX6124);
	not 	XG11688 	(WX6123,WX6122);
	not 	XG11689 	(WX6121,WX6120);
	not 	XG11690 	(WX6119,WX6118);
	not 	XG11691 	(WX6117,WX6116);
	not 	XG11692 	(WX6115,WX6114);
	not 	XG11693 	(WX6113,WX6112);
	not 	XG11694 	(WX6111,WX6110);
	not 	XG11695 	(WX6109,WX6108);
	not 	XG11696 	(WX6107,WX6106);
	not 	XG11697 	(WX6105,WX6104);
	not 	XG11698 	(WX6167,WX6166);
	not 	XG11699 	(WX6165,WX6164);
	not 	XG11700 	(WX6163,WX6162);
	not 	XG11701 	(WX6161,WX6160);
	not 	XG11702 	(WX6159,WX6158);
	not 	XG11703 	(WX6157,WX6156);
	not 	XG11704 	(WX6155,WX6154);
	not 	XG11705 	(WX6153,WX6152);
	not 	XG11706 	(WX6151,WX6150);
	not 	XG11707 	(WX6149,WX6148);
	not 	XG11708 	(WX6147,WX6146);
	not 	XG11709 	(WX6145,WX6144);
	not 	XG11710 	(WX6143,WX6142);
	not 	XG11711 	(WX6141,WX6140);
	not 	XG11712 	(WX6139,WX6138);
	not 	XG11713 	(WX6137,WX6136);
	not 	XG11714 	(WX4842,WX4841);
	not 	XG11715 	(WX4840,WX4839);
	not 	XG11716 	(WX4838,WX4837);
	not 	XG11717 	(WX4836,WX4835);
	not 	XG11718 	(WX4834,WX4833);
	not 	XG11719 	(WX4832,WX4831);
	not 	XG11720 	(WX4830,WX4829);
	not 	XG11721 	(WX4828,WX4827);
	not 	XG11722 	(WX4826,WX4825);
	not 	XG11723 	(WX4824,WX4823);
	not 	XG11724 	(WX4822,WX4821);
	not 	XG11725 	(WX4820,WX4819);
	not 	XG11726 	(WX4818,WX4817);
	not 	XG11727 	(WX4816,WX4815);
	not 	XG11728 	(WX4814,WX4813);
	not 	XG11729 	(WX4812,WX4811);
	not 	XG11730 	(WX4874,WX4873);
	not 	XG11731 	(WX4872,WX4871);
	not 	XG11732 	(WX4870,WX4869);
	not 	XG11733 	(WX4868,WX4867);
	not 	XG11734 	(WX4866,WX4865);
	not 	XG11735 	(WX4864,WX4863);
	not 	XG11736 	(WX4862,WX4861);
	not 	XG11737 	(WX4860,WX4859);
	not 	XG11738 	(WX4858,WX4857);
	not 	XG11739 	(WX4856,WX4855);
	not 	XG11740 	(WX4854,WX4853);
	not 	XG11741 	(WX4852,WX4851);
	not 	XG11742 	(WX4850,WX4849);
	not 	XG11743 	(WX4848,WX4847);
	not 	XG11744 	(WX4846,WX4845);
	not 	XG11745 	(WX4844,WX4843);
	not 	XG11746 	(WX3549,WX3548);
	not 	XG11747 	(WX3547,WX3546);
	not 	XG11748 	(WX3545,WX3544);
	not 	XG11749 	(WX3543,WX3542);
	not 	XG11750 	(WX3541,WX3540);
	not 	XG11751 	(WX3539,WX3538);
	not 	XG11752 	(WX3537,WX3536);
	not 	XG11753 	(WX3535,WX3534);
	not 	XG11754 	(WX3533,WX3532);
	not 	XG11755 	(WX3531,WX3530);
	not 	XG11756 	(WX3529,WX3528);
	not 	XG11757 	(WX3527,WX3526);
	not 	XG11758 	(WX3525,WX3524);
	not 	XG11759 	(WX3523,WX3522);
	not 	XG11760 	(WX3521,WX3520);
	not 	XG11761 	(WX3519,WX3518);
	not 	XG11762 	(WX3581,WX3580);
	not 	XG11763 	(WX3579,WX3578);
	not 	XG11764 	(WX3577,WX3576);
	not 	XG11765 	(WX3575,WX3574);
	not 	XG11766 	(WX3573,WX3572);
	not 	XG11767 	(WX3571,WX3570);
	not 	XG11768 	(WX3569,WX3568);
	not 	XG11769 	(WX3567,WX3566);
	not 	XG11770 	(WX3565,WX3564);
	not 	XG11771 	(WX3563,WX3562);
	not 	XG11772 	(WX3561,WX3560);
	not 	XG11773 	(WX3559,WX3558);
	not 	XG11774 	(WX3557,WX3556);
	not 	XG11775 	(WX3555,WX3554);
	not 	XG11776 	(WX3553,WX3552);
	not 	XG11777 	(WX3551,WX3550);
	not 	XG11778 	(WX2256,WX2255);
	not 	XG11779 	(WX2254,WX2253);
	not 	XG11780 	(WX2252,WX2251);
	not 	XG11781 	(WX2250,WX2249);
	not 	XG11782 	(WX2248,WX2247);
	not 	XG11783 	(WX2246,WX2245);
	not 	XG11784 	(WX2244,WX2243);
	not 	XG11785 	(WX2242,WX2241);
	not 	XG11786 	(WX2240,WX2239);
	not 	XG11787 	(WX2238,WX2237);
	not 	XG11788 	(WX2236,WX2235);
	not 	XG11789 	(WX2234,WX2233);
	not 	XG11790 	(WX2232,WX2231);
	not 	XG11791 	(WX2230,WX2229);
	not 	XG11792 	(WX2228,WX2227);
	not 	XG11793 	(WX2226,WX2225);
	not 	XG11794 	(WX2288,WX2287);
	not 	XG11795 	(WX2286,WX2285);
	not 	XG11796 	(WX2284,WX2283);
	not 	XG11797 	(WX2282,WX2281);
	not 	XG11798 	(WX2280,WX2279);
	not 	XG11799 	(WX2278,WX2277);
	not 	XG11800 	(WX2276,WX2275);
	not 	XG11801 	(WX2274,WX2273);
	not 	XG11802 	(WX2272,WX2271);
	not 	XG11803 	(WX2270,WX2269);
	not 	XG11804 	(WX2268,WX2267);
	not 	XG11805 	(WX2266,WX2265);
	not 	XG11806 	(WX2264,WX2263);
	not 	XG11807 	(WX2262,WX2261);
	not 	XG11808 	(WX2260,WX2259);
	not 	XG11809 	(WX2258,WX2257);
	not 	XG11810 	(WX963,WX962);
	not 	XG11811 	(WX961,WX960);
	not 	XG11812 	(WX959,WX958);
	not 	XG11813 	(WX957,WX956);
	not 	XG11814 	(WX955,WX954);
	not 	XG11815 	(WX953,WX952);
	not 	XG11816 	(WX951,WX950);
	not 	XG11817 	(WX949,WX948);
	not 	XG11818 	(WX947,WX946);
	not 	XG11819 	(WX945,WX944);
	not 	XG11820 	(WX943,WX942);
	not 	XG11821 	(WX941,WX940);
	not 	XG11822 	(WX939,WX938);
	not 	XG11823 	(WX937,WX936);
	not 	XG11824 	(WX935,WX934);
	not 	XG11825 	(WX933,WX932);
	not 	XG11826 	(WX995,WX994);
	not 	XG11827 	(WX993,WX992);
	not 	XG11828 	(WX991,WX990);
	not 	XG11829 	(WX989,WX988);
	not 	XG11830 	(WX987,WX986);
	not 	XG11831 	(WX985,WX984);
	not 	XG11832 	(WX983,WX982);
	not 	XG11833 	(WX981,WX980);
	not 	XG11834 	(WX979,WX978);
	not 	XG11835 	(WX977,WX976);
	not 	XG11836 	(WX975,WX974);
	not 	XG11837 	(WX973,WX972);
	not 	XG11838 	(WX971,WX970);
	not 	XG11839 	(WX969,WX968);
	not 	XG11840 	(WX967,WX966);
	not 	XG11841 	(WX965,WX964);
	not 	XG11842 	(WX548,WX965);
	not 	XG11843 	(WX549,WX967);
	not 	XG11844 	(WX550,WX969);
	not 	XG11845 	(WX551,WX971);
	not 	XG11846 	(WX552,WX973);
	not 	XG11847 	(WX553,WX975);
	not 	XG11848 	(WX554,WX977);
	not 	XG11849 	(WX555,WX979);
	not 	XG11850 	(WX556,WX981);
	not 	XG11851 	(WX557,WX983);
	not 	XG11852 	(WX558,WX985);
	not 	XG11853 	(WX559,WX987);
	not 	XG11854 	(WX560,WX989);
	not 	XG11855 	(WX561,WX991);
	not 	XG11856 	(WX562,WX993);
	not 	XG11857 	(WX563,WX995);
	not 	XG11858 	(WX564,WX933);
	not 	XG11859 	(WX565,WX935);
	not 	XG11860 	(WX566,WX937);
	not 	XG11861 	(WX567,WX939);
	not 	XG11862 	(WX568,WX941);
	not 	XG11863 	(WX569,WX943);
	not 	XG11864 	(WX570,WX945);
	not 	XG11865 	(WX571,WX947);
	not 	XG11866 	(WX572,WX949);
	not 	XG11867 	(WX573,WX951);
	not 	XG11868 	(WX574,WX953);
	not 	XG11869 	(WX575,WX955);
	not 	XG11870 	(WX576,WX957);
	not 	XG11871 	(WX577,WX959);
	not 	XG11872 	(WX578,WX961);
	not 	XG11873 	(WX579,WX963);
	not 	XG11874 	(WX1841,WX2258);
	not 	XG11875 	(WX1842,WX2260);
	not 	XG11876 	(WX1843,WX2262);
	not 	XG11877 	(WX1844,WX2264);
	not 	XG11878 	(WX1845,WX2266);
	not 	XG11879 	(WX1846,WX2268);
	not 	XG11880 	(WX1847,WX2270);
	not 	XG11881 	(WX1848,WX2272);
	not 	XG11882 	(WX1849,WX2274);
	not 	XG11883 	(WX1850,WX2276);
	not 	XG11884 	(WX1851,WX2278);
	not 	XG11885 	(WX1852,WX2280);
	not 	XG11886 	(WX1853,WX2282);
	not 	XG11887 	(WX1854,WX2284);
	not 	XG11888 	(WX1855,WX2286);
	not 	XG11889 	(WX1856,WX2288);
	not 	XG11890 	(WX1857,WX2226);
	not 	XG11891 	(WX1858,WX2228);
	not 	XG11892 	(WX1859,WX2230);
	not 	XG11893 	(WX1860,WX2232);
	not 	XG11894 	(WX1861,WX2234);
	not 	XG11895 	(WX1862,WX2236);
	not 	XG11896 	(WX1863,WX2238);
	not 	XG11897 	(WX1864,WX2240);
	not 	XG11898 	(WX1865,WX2242);
	not 	XG11899 	(WX1866,WX2244);
	not 	XG11900 	(WX1867,WX2246);
	not 	XG11901 	(WX1868,WX2248);
	not 	XG11902 	(WX1869,WX2250);
	not 	XG11903 	(WX1870,WX2252);
	not 	XG11904 	(WX1871,WX2254);
	not 	XG11905 	(WX1872,WX2256);
	not 	XG11906 	(WX3134,WX3551);
	not 	XG11907 	(WX3135,WX3553);
	not 	XG11908 	(WX3136,WX3555);
	not 	XG11909 	(WX3137,WX3557);
	not 	XG11910 	(WX3138,WX3559);
	not 	XG11911 	(WX3139,WX3561);
	not 	XG11912 	(WX3140,WX3563);
	not 	XG11913 	(WX3141,WX3565);
	not 	XG11914 	(WX3142,WX3567);
	not 	XG11915 	(WX3143,WX3569);
	not 	XG11916 	(WX3144,WX3571);
	not 	XG11917 	(WX3145,WX3573);
	not 	XG11918 	(WX3146,WX3575);
	not 	XG11919 	(WX3147,WX3577);
	not 	XG11920 	(WX3148,WX3579);
	not 	XG11921 	(WX3149,WX3581);
	not 	XG11922 	(WX3150,WX3519);
	not 	XG11923 	(WX3151,WX3521);
	not 	XG11924 	(WX3152,WX3523);
	not 	XG11925 	(WX3153,WX3525);
	not 	XG11926 	(WX3154,WX3527);
	not 	XG11927 	(WX3155,WX3529);
	not 	XG11928 	(WX3156,WX3531);
	not 	XG11929 	(WX3157,WX3533);
	not 	XG11930 	(WX3158,WX3535);
	not 	XG11931 	(WX3159,WX3537);
	not 	XG11932 	(WX3160,WX3539);
	not 	XG11933 	(WX3161,WX3541);
	not 	XG11934 	(WX3162,WX3543);
	not 	XG11935 	(WX3163,WX3545);
	not 	XG11936 	(WX3164,WX3547);
	not 	XG11937 	(WX3165,WX3549);
	not 	XG11938 	(WX4427,WX4844);
	not 	XG11939 	(WX4428,WX4846);
	not 	XG11940 	(WX4429,WX4848);
	not 	XG11941 	(WX4430,WX4850);
	not 	XG11942 	(WX4431,WX4852);
	not 	XG11943 	(WX4432,WX4854);
	not 	XG11944 	(WX4433,WX4856);
	not 	XG11945 	(WX4434,WX4858);
	not 	XG11946 	(WX4435,WX4860);
	not 	XG11947 	(WX4436,WX4862);
	not 	XG11948 	(WX4437,WX4864);
	not 	XG11949 	(WX4438,WX4866);
	not 	XG11950 	(WX4439,WX4868);
	not 	XG11951 	(WX4440,WX4870);
	not 	XG11952 	(WX4441,WX4872);
	not 	XG11953 	(WX4442,WX4874);
	not 	XG11954 	(WX4443,WX4812);
	not 	XG11955 	(WX4444,WX4814);
	not 	XG11956 	(WX4445,WX4816);
	not 	XG11957 	(WX4446,WX4818);
	not 	XG11958 	(WX4447,WX4820);
	not 	XG11959 	(WX4448,WX4822);
	not 	XG11960 	(WX4449,WX4824);
	not 	XG11961 	(WX4450,WX4826);
	not 	XG11962 	(WX4451,WX4828);
	not 	XG11963 	(WX4452,WX4830);
	not 	XG11964 	(WX4453,WX4832);
	not 	XG11965 	(WX4454,WX4834);
	not 	XG11966 	(WX4455,WX4836);
	not 	XG11967 	(WX4456,WX4838);
	not 	XG11968 	(WX4457,WX4840);
	not 	XG11969 	(WX4458,WX4842);
	not 	XG11970 	(WX5720,WX6137);
	not 	XG11971 	(WX5721,WX6139);
	not 	XG11972 	(WX5722,WX6141);
	not 	XG11973 	(WX5723,WX6143);
	not 	XG11974 	(WX5724,WX6145);
	not 	XG11975 	(WX5725,WX6147);
	not 	XG11976 	(WX5726,WX6149);
	not 	XG11977 	(WX5727,WX6151);
	not 	XG11978 	(WX5728,WX6153);
	not 	XG11979 	(WX5729,WX6155);
	not 	XG11980 	(WX5730,WX6157);
	not 	XG11981 	(WX5731,WX6159);
	not 	XG11982 	(WX5732,WX6161);
	not 	XG11983 	(WX5733,WX6163);
	not 	XG11984 	(WX5734,WX6165);
	not 	XG11985 	(WX5735,WX6167);
	not 	XG11986 	(WX5736,WX6105);
	not 	XG11987 	(WX5737,WX6107);
	not 	XG11988 	(WX5738,WX6109);
	not 	XG11989 	(WX5739,WX6111);
	not 	XG11990 	(WX5740,WX6113);
	not 	XG11991 	(WX5741,WX6115);
	not 	XG11992 	(WX5742,WX6117);
	not 	XG11993 	(WX5743,WX6119);
	not 	XG11994 	(WX5744,WX6121);
	not 	XG11995 	(WX5745,WX6123);
	not 	XG11996 	(WX5746,WX6125);
	not 	XG11997 	(WX5747,WX6127);
	not 	XG11998 	(WX5748,WX6129);
	not 	XG11999 	(WX5749,WX6131);
	not 	XG12000 	(WX5750,WX6133);
	not 	XG12001 	(WX5751,WX6135);
	not 	XG12002 	(WX7013,WX7430);
	not 	XG12003 	(WX7014,WX7432);
	not 	XG12004 	(WX7015,WX7434);
	not 	XG12005 	(WX7016,WX7436);
	not 	XG12006 	(WX7017,WX7438);
	not 	XG12007 	(WX7018,WX7440);
	not 	XG12008 	(WX7019,WX7442);
	not 	XG12009 	(WX7020,WX7444);
	not 	XG12010 	(WX7021,WX7446);
	not 	XG12011 	(WX7022,WX7448);
	not 	XG12012 	(WX7023,WX7450);
	not 	XG12013 	(WX7024,WX7452);
	not 	XG12014 	(WX7025,WX7454);
	not 	XG12015 	(WX7026,WX7456);
	not 	XG12016 	(WX7027,WX7458);
	not 	XG12017 	(WX7028,WX7460);
	not 	XG12018 	(WX7029,WX7398);
	not 	XG12019 	(WX7030,WX7400);
	not 	XG12020 	(WX7031,WX7402);
	not 	XG12021 	(WX7032,WX7404);
	not 	XG12022 	(WX7033,WX7406);
	not 	XG12023 	(WX7034,WX7408);
	not 	XG12024 	(WX7035,WX7410);
	not 	XG12025 	(WX7036,WX7412);
	not 	XG12026 	(WX7037,WX7414);
	not 	XG12027 	(WX7038,WX7416);
	not 	XG12028 	(WX7039,WX7418);
	not 	XG12029 	(WX7040,WX7420);
	not 	XG12030 	(WX7041,WX7422);
	not 	XG12031 	(WX7042,WX7424);
	not 	XG12032 	(WX7043,WX7426);
	not 	XG12033 	(WX7044,WX7428);
	not 	XG12034 	(WX8306,WX8723);
	not 	XG12035 	(WX8307,WX8725);
	not 	XG12036 	(WX8308,WX8727);
	not 	XG12037 	(WX8309,WX8729);
	not 	XG12038 	(WX8310,WX8731);
	not 	XG12039 	(WX8311,WX8733);
	not 	XG12040 	(WX8312,WX8735);
	not 	XG12041 	(WX8313,WX8737);
	not 	XG12042 	(WX8314,WX8739);
	not 	XG12043 	(WX8315,WX8741);
	not 	XG12044 	(WX8316,WX8743);
	not 	XG12045 	(WX8317,WX8745);
	not 	XG12046 	(WX8318,WX8747);
	not 	XG12047 	(WX8319,WX8749);
	not 	XG12048 	(WX8320,WX8751);
	not 	XG12049 	(WX8321,WX8753);
	not 	XG12050 	(WX8322,WX8691);
	not 	XG12051 	(WX8323,WX8693);
	not 	XG12052 	(WX8324,WX8695);
	not 	XG12053 	(WX8325,WX8697);
	not 	XG12054 	(WX8326,WX8699);
	not 	XG12055 	(WX8327,WX8701);
	not 	XG12056 	(WX8328,WX8703);
	not 	XG12057 	(WX8329,WX8705);
	not 	XG12058 	(WX8330,WX8707);
	not 	XG12059 	(WX8331,WX8709);
	not 	XG12060 	(WX8332,WX8711);
	not 	XG12061 	(WX8333,WX8713);
	not 	XG12062 	(WX8334,WX8715);
	not 	XG12063 	(WX8335,WX8717);
	not 	XG12064 	(WX8336,WX8719);
	not 	XG12065 	(WX8337,WX8721);
	not 	XG12066 	(WX9599,WX10016);
	not 	XG12067 	(WX9600,WX10018);
	not 	XG12068 	(WX9601,WX10020);
	not 	XG12069 	(WX9602,WX10022);
	not 	XG12070 	(WX9603,WX10024);
	not 	XG12071 	(WX9604,WX10026);
	not 	XG12072 	(WX9605,WX10028);
	not 	XG12073 	(WX9606,WX10030);
	not 	XG12074 	(WX9607,WX10032);
	not 	XG12075 	(WX9608,WX10034);
	not 	XG12076 	(WX9609,WX10036);
	not 	XG12077 	(WX9610,WX10038);
	not 	XG12078 	(WX9611,WX10040);
	not 	XG12079 	(WX9612,WX10042);
	not 	XG12080 	(WX9613,WX10044);
	not 	XG12081 	(WX9614,WX10046);
	not 	XG12082 	(WX9615,WX9984);
	not 	XG12083 	(WX9616,WX9986);
	not 	XG12084 	(WX9617,WX9988);
	not 	XG12085 	(WX9618,WX9990);
	not 	XG12086 	(WX9619,WX9992);
	not 	XG12087 	(WX9620,WX9994);
	not 	XG12088 	(WX9621,WX9996);
	not 	XG12089 	(WX9622,WX9998);
	not 	XG12090 	(WX9623,WX10000);
	not 	XG12091 	(WX9624,WX10002);
	not 	XG12092 	(WX9625,WX10004);
	not 	XG12093 	(WX9626,WX10006);
	not 	XG12094 	(WX9627,WX10008);
	not 	XG12095 	(WX9628,WX10010);
	not 	XG12096 	(WX9629,WX10012);
	not 	XG12097 	(WX9630,WX10014);
	not 	XG12098 	(WX10892,WX11309);
	not 	XG12099 	(WX10893,WX11311);
	not 	XG12100 	(WX10894,WX11313);
	not 	XG12101 	(WX10895,WX11315);
	not 	XG12102 	(WX10896,WX11317);
	not 	XG12103 	(WX10897,WX11319);
	not 	XG12104 	(WX10898,WX11321);
	not 	XG12105 	(WX10899,WX11323);
	not 	XG12106 	(WX10900,WX11325);
	not 	XG12107 	(WX10901,WX11327);
	not 	XG12108 	(WX10902,WX11329);
	not 	XG12109 	(WX10903,WX11331);
	not 	XG12110 	(WX10904,WX11333);
	not 	XG12111 	(WX10905,WX11335);
	not 	XG12112 	(WX10906,WX11337);
	not 	XG12113 	(WX10907,WX11339);
	not 	XG12114 	(WX10908,WX11277);
	not 	XG12115 	(WX10909,WX11279);
	not 	XG12116 	(WX10910,WX11281);
	not 	XG12117 	(WX10911,WX11283);
	not 	XG12118 	(WX10912,WX11285);
	not 	XG12119 	(WX10913,WX11287);
	not 	XG12120 	(WX10914,WX11289);
	not 	XG12121 	(WX10915,WX11291);
	not 	XG12122 	(WX10916,WX11293);
	not 	XG12123 	(WX10917,WX11295);
	not 	XG12124 	(WX10918,WX11297);
	not 	XG12125 	(WX10919,WX11299);
	not 	XG12126 	(WX10920,WX11301);
	not 	XG12127 	(WX10921,WX11303);
	not 	XG12128 	(WX10922,WX11305);
	not 	XG12129 	(WX10923,WX11307);
	not 	XG12130 	(WX10955,WX10923);
	not 	XG12131 	(WX10954,WX10922);
	not 	XG12132 	(WX10953,WX10921);
	not 	XG12133 	(WX10952,WX10920);
	not 	XG12134 	(WX10951,WX10919);
	not 	XG12135 	(WX10950,WX10918);
	not 	XG12136 	(WX10949,WX10917);
	not 	XG12137 	(WX10948,WX10916);
	not 	XG12138 	(WX10947,WX10915);
	not 	XG12139 	(WX10946,WX10914);
	not 	XG12140 	(WX10945,WX10913);
	not 	XG12141 	(WX10944,WX10912);
	not 	XG12142 	(WX10943,WX10911);
	not 	XG12143 	(WX10942,WX10910);
	not 	XG12144 	(WX10941,WX10909);
	not 	XG12145 	(WX10940,WX10908);
	not 	XG12146 	(WX10939,WX10907);
	not 	XG12147 	(WX10938,WX10906);
	not 	XG12148 	(WX10937,WX10905);
	not 	XG12149 	(WX10936,WX10904);
	not 	XG12150 	(WX10935,WX10903);
	not 	XG12151 	(WX10934,WX10902);
	not 	XG12152 	(WX10933,WX10901);
	not 	XG12153 	(WX10932,WX10900);
	not 	XG12154 	(WX10931,WX10899);
	not 	XG12155 	(WX10930,WX10898);
	not 	XG12156 	(WX10929,WX10897);
	not 	XG12157 	(WX10928,WX10896);
	not 	XG12158 	(WX10927,WX10895);
	not 	XG12159 	(WX10926,WX10894);
	not 	XG12160 	(WX10925,WX10893);
	not 	XG12161 	(WX10924,WX10892);
	not 	XG12162 	(WX9662,WX9630);
	not 	XG12163 	(WX9661,WX9629);
	not 	XG12164 	(WX9660,WX9628);
	not 	XG12165 	(WX9659,WX9627);
	not 	XG12166 	(WX9658,WX9626);
	not 	XG12167 	(WX9657,WX9625);
	not 	XG12168 	(WX9656,WX9624);
	not 	XG12169 	(WX9655,WX9623);
	not 	XG12170 	(WX9654,WX9622);
	not 	XG12171 	(WX9653,WX9621);
	not 	XG12172 	(WX9652,WX9620);
	not 	XG12173 	(WX9651,WX9619);
	not 	XG12174 	(WX9650,WX9618);
	not 	XG12175 	(WX9649,WX9617);
	not 	XG12176 	(WX9648,WX9616);
	not 	XG12177 	(WX9647,WX9615);
	not 	XG12178 	(WX9646,WX9614);
	not 	XG12179 	(WX9645,WX9613);
	not 	XG12180 	(WX9644,WX9612);
	not 	XG12181 	(WX9643,WX9611);
	not 	XG12182 	(WX9642,WX9610);
	not 	XG12183 	(WX9641,WX9609);
	not 	XG12184 	(WX9640,WX9608);
	not 	XG12185 	(WX9639,WX9607);
	not 	XG12186 	(WX9638,WX9606);
	not 	XG12187 	(WX9637,WX9605);
	not 	XG12188 	(WX9636,WX9604);
	not 	XG12189 	(WX9635,WX9603);
	not 	XG12190 	(WX9634,WX9602);
	not 	XG12191 	(WX9633,WX9601);
	not 	XG12192 	(WX9632,WX9600);
	not 	XG12193 	(WX9631,WX9599);
	not 	XG12194 	(WX8369,WX8337);
	not 	XG12195 	(WX8368,WX8336);
	not 	XG12196 	(WX8367,WX8335);
	not 	XG12197 	(WX8366,WX8334);
	not 	XG12198 	(WX8365,WX8333);
	not 	XG12199 	(WX8364,WX8332);
	not 	XG12200 	(WX8363,WX8331);
	not 	XG12201 	(WX8362,WX8330);
	not 	XG12202 	(WX8361,WX8329);
	not 	XG12203 	(WX8360,WX8328);
	not 	XG12204 	(WX8359,WX8327);
	not 	XG12205 	(WX8358,WX8326);
	not 	XG12206 	(WX8357,WX8325);
	not 	XG12207 	(WX8356,WX8324);
	not 	XG12208 	(WX8355,WX8323);
	not 	XG12209 	(WX8354,WX8322);
	not 	XG12210 	(WX8353,WX8321);
	not 	XG12211 	(WX8352,WX8320);
	not 	XG12212 	(WX8351,WX8319);
	not 	XG12213 	(WX8350,WX8318);
	not 	XG12214 	(WX8349,WX8317);
	not 	XG12215 	(WX8348,WX8316);
	not 	XG12216 	(WX8347,WX8315);
	not 	XG12217 	(WX8346,WX8314);
	not 	XG12218 	(WX8345,WX8313);
	not 	XG12219 	(WX8344,WX8312);
	not 	XG12220 	(WX8343,WX8311);
	not 	XG12221 	(WX8342,WX8310);
	not 	XG12222 	(WX8341,WX8309);
	not 	XG12223 	(WX8340,WX8308);
	not 	XG12224 	(WX8339,WX8307);
	not 	XG12225 	(WX8338,WX8306);
	not 	XG12226 	(WX7076,WX7044);
	not 	XG12227 	(WX7075,WX7043);
	not 	XG12228 	(WX7074,WX7042);
	not 	XG12229 	(WX7073,WX7041);
	not 	XG12230 	(WX7072,WX7040);
	not 	XG12231 	(WX7071,WX7039);
	not 	XG12232 	(WX7070,WX7038);
	not 	XG12233 	(WX7069,WX7037);
	not 	XG12234 	(WX7068,WX7036);
	not 	XG12235 	(WX7067,WX7035);
	not 	XG12236 	(WX7066,WX7034);
	not 	XG12237 	(WX7065,WX7033);
	not 	XG12238 	(WX7064,WX7032);
	not 	XG12239 	(WX7063,WX7031);
	not 	XG12240 	(WX7062,WX7030);
	not 	XG12241 	(WX7061,WX7029);
	not 	XG12242 	(WX7060,WX7028);
	not 	XG12243 	(WX7059,WX7027);
	not 	XG12244 	(WX7058,WX7026);
	not 	XG12245 	(WX7057,WX7025);
	not 	XG12246 	(WX7056,WX7024);
	not 	XG12247 	(WX7055,WX7023);
	not 	XG12248 	(WX7054,WX7022);
	not 	XG12249 	(WX7053,WX7021);
	not 	XG12250 	(WX7052,WX7020);
	not 	XG12251 	(WX7051,WX7019);
	not 	XG12252 	(WX7050,WX7018);
	not 	XG12253 	(WX7049,WX7017);
	not 	XG12254 	(WX7048,WX7016);
	not 	XG12255 	(WX7047,WX7015);
	not 	XG12256 	(WX7046,WX7014);
	not 	XG12257 	(WX7045,WX7013);
	not 	XG12258 	(WX5783,WX5751);
	not 	XG12259 	(WX5782,WX5750);
	not 	XG12260 	(WX5781,WX5749);
	not 	XG12261 	(WX5780,WX5748);
	not 	XG12262 	(WX5779,WX5747);
	not 	XG12263 	(WX5778,WX5746);
	not 	XG12264 	(WX5777,WX5745);
	not 	XG12265 	(WX5776,WX5744);
	not 	XG12266 	(WX5775,WX5743);
	not 	XG12267 	(WX5774,WX5742);
	not 	XG12268 	(WX5773,WX5741);
	not 	XG12269 	(WX5772,WX5740);
	not 	XG12270 	(WX5771,WX5739);
	not 	XG12271 	(WX5770,WX5738);
	not 	XG12272 	(WX5769,WX5737);
	not 	XG12273 	(WX5768,WX5736);
	not 	XG12274 	(WX5767,WX5735);
	not 	XG12275 	(WX5766,WX5734);
	not 	XG12276 	(WX5765,WX5733);
	not 	XG12277 	(WX5764,WX5732);
	not 	XG12278 	(WX5763,WX5731);
	not 	XG12279 	(WX5762,WX5730);
	not 	XG12280 	(WX5761,WX5729);
	not 	XG12281 	(WX5760,WX5728);
	not 	XG12282 	(WX5759,WX5727);
	not 	XG12283 	(WX5758,WX5726);
	not 	XG12284 	(WX5757,WX5725);
	not 	XG12285 	(WX5756,WX5724);
	not 	XG12286 	(WX5755,WX5723);
	not 	XG12287 	(WX5754,WX5722);
	not 	XG12288 	(WX5753,WX5721);
	not 	XG12289 	(WX5752,WX5720);
	not 	XG12290 	(WX4490,WX4458);
	not 	XG12291 	(WX4489,WX4457);
	not 	XG12292 	(WX4488,WX4456);
	not 	XG12293 	(WX4487,WX4455);
	not 	XG12294 	(WX4486,WX4454);
	not 	XG12295 	(WX4485,WX4453);
	not 	XG12296 	(WX4484,WX4452);
	not 	XG12297 	(WX4483,WX4451);
	not 	XG12298 	(WX4482,WX4450);
	not 	XG12299 	(WX4481,WX4449);
	not 	XG12300 	(WX4480,WX4448);
	not 	XG12301 	(WX4479,WX4447);
	not 	XG12302 	(WX4478,WX4446);
	not 	XG12303 	(WX4477,WX4445);
	not 	XG12304 	(WX4476,WX4444);
	not 	XG12305 	(WX4475,WX4443);
	not 	XG12306 	(WX4474,WX4442);
	not 	XG12307 	(WX4473,WX4441);
	not 	XG12308 	(WX4472,WX4440);
	not 	XG12309 	(WX4471,WX4439);
	not 	XG12310 	(WX4470,WX4438);
	not 	XG12311 	(WX4469,WX4437);
	not 	XG12312 	(WX4468,WX4436);
	not 	XG12313 	(WX4467,WX4435);
	not 	XG12314 	(WX4466,WX4434);
	not 	XG12315 	(WX4465,WX4433);
	not 	XG12316 	(WX4464,WX4432);
	not 	XG12317 	(WX4463,WX4431);
	not 	XG12318 	(WX4462,WX4430);
	not 	XG12319 	(WX4461,WX4429);
	not 	XG12320 	(WX4460,WX4428);
	not 	XG12321 	(WX4459,WX4427);
	not 	XG12322 	(WX3197,WX3165);
	not 	XG12323 	(WX3196,WX3164);
	not 	XG12324 	(WX3195,WX3163);
	not 	XG12325 	(WX3194,WX3162);
	not 	XG12326 	(WX3193,WX3161);
	not 	XG12327 	(WX3192,WX3160);
	not 	XG12328 	(WX3191,WX3159);
	not 	XG12329 	(WX3190,WX3158);
	not 	XG12330 	(WX3189,WX3157);
	not 	XG12331 	(WX3188,WX3156);
	not 	XG12332 	(WX3187,WX3155);
	not 	XG12333 	(WX3186,WX3154);
	not 	XG12334 	(WX3185,WX3153);
	not 	XG12335 	(WX3184,WX3152);
	not 	XG12336 	(WX3183,WX3151);
	not 	XG12337 	(WX3182,WX3150);
	not 	XG12338 	(WX3181,WX3149);
	not 	XG12339 	(WX3180,WX3148);
	not 	XG12340 	(WX3179,WX3147);
	not 	XG12341 	(WX3178,WX3146);
	not 	XG12342 	(WX3177,WX3145);
	not 	XG12343 	(WX3176,WX3144);
	not 	XG12344 	(WX3175,WX3143);
	not 	XG12345 	(WX3174,WX3142);
	not 	XG12346 	(WX3173,WX3141);
	not 	XG12347 	(WX3172,WX3140);
	not 	XG12348 	(WX3171,WX3139);
	not 	XG12349 	(WX3170,WX3138);
	not 	XG12350 	(WX3169,WX3137);
	not 	XG12351 	(WX3168,WX3136);
	not 	XG12352 	(WX3167,WX3135);
	not 	XG12353 	(WX3166,WX3134);
	not 	XG12354 	(WX1904,WX1872);
	not 	XG12355 	(WX1903,WX1871);
	not 	XG12356 	(WX1902,WX1870);
	not 	XG12357 	(WX1901,WX1869);
	not 	XG12358 	(WX1900,WX1868);
	not 	XG12359 	(WX1899,WX1867);
	not 	XG12360 	(WX1898,WX1866);
	not 	XG12361 	(WX1897,WX1865);
	not 	XG12362 	(WX1896,WX1864);
	not 	XG12363 	(WX1895,WX1863);
	not 	XG12364 	(WX1894,WX1862);
	not 	XG12365 	(WX1893,WX1861);
	not 	XG12366 	(WX1892,WX1860);
	not 	XG12367 	(WX1891,WX1859);
	not 	XG12368 	(WX1890,WX1858);
	not 	XG12369 	(WX1889,WX1857);
	not 	XG12370 	(WX1888,WX1856);
	not 	XG12371 	(WX1887,WX1855);
	not 	XG12372 	(WX1886,WX1854);
	not 	XG12373 	(WX1885,WX1853);
	not 	XG12374 	(WX1884,WX1852);
	not 	XG12375 	(WX1883,WX1851);
	not 	XG12376 	(WX1882,WX1850);
	not 	XG12377 	(WX1881,WX1849);
	not 	XG12378 	(WX1880,WX1848);
	not 	XG12379 	(WX1879,WX1847);
	not 	XG12380 	(WX1878,WX1846);
	not 	XG12381 	(WX1877,WX1845);
	not 	XG12382 	(WX1876,WX1844);
	not 	XG12383 	(WX1875,WX1843);
	not 	XG12384 	(WX1874,WX1842);
	not 	XG12385 	(WX1873,WX1841);
	not 	XG12386 	(WX611,WX579);
	not 	XG12387 	(WX610,WX578);
	not 	XG12388 	(WX609,WX577);
	not 	XG12389 	(WX608,WX576);
	not 	XG12390 	(WX607,WX575);
	not 	XG12391 	(WX606,WX574);
	not 	XG12392 	(WX605,WX573);
	not 	XG12393 	(WX604,WX572);
	not 	XG12394 	(WX603,WX571);
	not 	XG12395 	(WX602,WX570);
	not 	XG12396 	(WX601,WX569);
	not 	XG12397 	(WX600,WX568);
	not 	XG12398 	(WX599,WX567);
	not 	XG12399 	(WX598,WX566);
	not 	XG12400 	(WX597,WX565);
	not 	XG12401 	(WX596,WX564);
	not 	XG12402 	(WX595,WX563);
	not 	XG12403 	(WX594,WX562);
	not 	XG12404 	(WX593,WX561);
	not 	XG12405 	(WX592,WX560);
	not 	XG12406 	(WX591,WX559);
	not 	XG12407 	(WX590,WX558);
	not 	XG12408 	(WX589,WX557);
	not 	XG12409 	(WX588,WX556);
	not 	XG12410 	(WX587,WX555);
	not 	XG12411 	(WX586,WX554);
	not 	XG12412 	(WX585,WX553);
	not 	XG12413 	(WX584,WX552);
	not 	XG12414 	(WX583,WX551);
	not 	XG12415 	(WX582,WX550);
	not 	XG12416 	(WX581,WX549);
	not 	XG12417 	(WX580,WX548);
	and 	XG12418 	(WX11569,WX11570,WX10955);
	and 	XG12419 	(WX11562,WX11563,WX10954);
	and 	XG12420 	(WX11555,WX11556,WX10953);
	and 	XG12421 	(WX11548,WX11549,WX10952);
	and 	XG12422 	(WX11541,WX11542,WX10951);
	and 	XG12423 	(WX11534,WX11535,WX10950);
	and 	XG12424 	(WX11527,WX11528,WX10949);
	and 	XG12425 	(WX11520,WX11521,WX10948);
	and 	XG12426 	(WX11513,WX11514,WX10947);
	and 	XG12427 	(WX11506,WX11507,WX10946);
	and 	XG12428 	(WX11499,WX11500,WX10945);
	and 	XG12429 	(WX11492,WX11493,WX10944);
	and 	XG12430 	(WX11485,WX11486,WX10943);
	and 	XG12431 	(WX11478,WX11479,WX10942);
	and 	XG12432 	(WX11471,WX11472,WX10941);
	and 	XG12433 	(WX11464,WX11465,WX10940);
	and 	XG12434 	(WX11457,WX11458,WX10939);
	and 	XG12435 	(WX11450,WX11451,WX10938);
	and 	XG12436 	(WX11443,WX11444,WX10937);
	and 	XG12437 	(WX11436,WX11437,WX10936);
	and 	XG12438 	(WX11429,WX11430,WX10935);
	and 	XG12439 	(WX11422,WX11423,WX10934);
	and 	XG12440 	(WX11415,WX11416,WX10933);
	and 	XG12441 	(WX11408,WX11409,WX10932);
	and 	XG12442 	(WX11401,WX11402,WX10931);
	and 	XG12443 	(WX11394,WX11395,WX10930);
	and 	XG12444 	(WX11387,WX11388,WX10929);
	and 	XG12445 	(WX11380,WX11381,WX10928);
	and 	XG12446 	(WX11373,WX11374,WX10927);
	and 	XG12447 	(WX11366,WX11367,WX10926);
	and 	XG12448 	(WX11359,WX11360,WX10925);
	and 	XG12449 	(WX11352,WX11353,WX10924);
	and 	XG12450 	(WX10276,WX10277,WX9662);
	and 	XG12451 	(WX10269,WX10270,WX9661);
	and 	XG12452 	(WX10262,WX10263,WX9660);
	and 	XG12453 	(WX10255,WX10256,WX9659);
	and 	XG12454 	(WX10248,WX10249,WX9658);
	and 	XG12455 	(WX10241,WX10242,WX9657);
	and 	XG12456 	(WX10234,WX10235,WX9656);
	and 	XG12457 	(WX10227,WX10228,WX9655);
	and 	XG12458 	(WX10220,WX10221,WX9654);
	and 	XG12459 	(WX10213,WX10214,WX9653);
	and 	XG12460 	(WX10206,WX10207,WX9652);
	and 	XG12461 	(WX10199,WX10200,WX9651);
	and 	XG12462 	(WX10192,WX10193,WX9650);
	and 	XG12463 	(WX10185,WX10186,WX9649);
	and 	XG12464 	(WX10178,WX10179,WX9648);
	and 	XG12465 	(WX10171,WX10172,WX9647);
	and 	XG12466 	(WX10164,WX10165,WX9646);
	and 	XG12467 	(WX10157,WX10158,WX9645);
	and 	XG12468 	(WX10150,WX10151,WX9644);
	and 	XG12469 	(WX10143,WX10144,WX9643);
	and 	XG12470 	(WX10136,WX10137,WX9642);
	and 	XG12471 	(WX10129,WX10130,WX9641);
	and 	XG12472 	(WX10122,WX10123,WX9640);
	and 	XG12473 	(WX10115,WX10116,WX9639);
	and 	XG12474 	(WX10108,WX10109,WX9638);
	and 	XG12475 	(WX10101,WX10102,WX9637);
	and 	XG12476 	(WX10094,WX10095,WX9636);
	and 	XG12477 	(WX10087,WX10088,WX9635);
	and 	XG12478 	(WX10080,WX10081,WX9634);
	and 	XG12479 	(WX10073,WX10074,WX9633);
	and 	XG12480 	(WX10066,WX10067,WX9632);
	and 	XG12481 	(WX10059,WX10060,WX9631);
	and 	XG12482 	(WX8983,WX8984,WX8369);
	and 	XG12483 	(WX8976,WX8977,WX8368);
	and 	XG12484 	(WX8969,WX8970,WX8367);
	and 	XG12485 	(WX8962,WX8963,WX8366);
	and 	XG12486 	(WX8955,WX8956,WX8365);
	and 	XG12487 	(WX8948,WX8949,WX8364);
	and 	XG12488 	(WX8941,WX8942,WX8363);
	and 	XG12489 	(WX8934,WX8935,WX8362);
	and 	XG12490 	(WX8927,WX8928,WX8361);
	and 	XG12491 	(WX8920,WX8921,WX8360);
	and 	XG12492 	(WX8913,WX8914,WX8359);
	and 	XG12493 	(WX8906,WX8907,WX8358);
	and 	XG12494 	(WX8899,WX8900,WX8357);
	and 	XG12495 	(WX8892,WX8893,WX8356);
	and 	XG12496 	(WX8885,WX8886,WX8355);
	and 	XG12497 	(WX8878,WX8879,WX8354);
	and 	XG12498 	(WX8871,WX8872,WX8353);
	and 	XG12499 	(WX8864,WX8865,WX8352);
	and 	XG12500 	(WX8857,WX8858,WX8351);
	and 	XG12501 	(WX8850,WX8851,WX8350);
	and 	XG12502 	(WX8843,WX8844,WX8349);
	and 	XG12503 	(WX8836,WX8837,WX8348);
	and 	XG12504 	(WX8829,WX8830,WX8347);
	and 	XG12505 	(WX8822,WX8823,WX8346);
	and 	XG12506 	(WX8815,WX8816,WX8345);
	and 	XG12507 	(WX8808,WX8809,WX8344);
	and 	XG12508 	(WX8801,WX8802,WX8343);
	and 	XG12509 	(WX8794,WX8795,WX8342);
	and 	XG12510 	(WX8787,WX8788,WX8341);
	and 	XG12511 	(WX8780,WX8781,WX8340);
	and 	XG12512 	(WX8773,WX8774,WX8339);
	and 	XG12513 	(WX8766,WX8767,WX8338);
	and 	XG12514 	(WX7690,WX7691,WX7076);
	and 	XG12515 	(WX7683,WX7684,WX7075);
	and 	XG12516 	(WX7676,WX7677,WX7074);
	and 	XG12517 	(WX7669,WX7670,WX7073);
	and 	XG12518 	(WX7662,WX7663,WX7072);
	and 	XG12519 	(WX7655,WX7656,WX7071);
	and 	XG12520 	(WX7648,WX7649,WX7070);
	and 	XG12521 	(WX7641,WX7642,WX7069);
	and 	XG12522 	(WX7634,WX7635,WX7068);
	and 	XG12523 	(WX7627,WX7628,WX7067);
	and 	XG12524 	(WX7620,WX7621,WX7066);
	and 	XG12525 	(WX7613,WX7614,WX7065);
	and 	XG12526 	(WX7606,WX7607,WX7064);
	and 	XG12527 	(WX7599,WX7600,WX7063);
	and 	XG12528 	(WX7592,WX7593,WX7062);
	and 	XG12529 	(WX7585,WX7586,WX7061);
	and 	XG12530 	(WX7578,WX7579,WX7060);
	and 	XG12531 	(WX7571,WX7572,WX7059);
	and 	XG12532 	(WX7564,WX7565,WX7058);
	and 	XG12533 	(WX7557,WX7558,WX7057);
	and 	XG12534 	(WX7550,WX7551,WX7056);
	and 	XG12535 	(WX7543,WX7544,WX7055);
	and 	XG12536 	(WX7536,WX7537,WX7054);
	and 	XG12537 	(WX7529,WX7530,WX7053);
	and 	XG12538 	(WX7522,WX7523,WX7052);
	and 	XG12539 	(WX7515,WX7516,WX7051);
	and 	XG12540 	(WX7508,WX7509,WX7050);
	and 	XG12541 	(WX7501,WX7502,WX7049);
	and 	XG12542 	(WX7494,WX7495,WX7048);
	and 	XG12543 	(WX7487,WX7488,WX7047);
	and 	XG12544 	(WX7480,WX7481,WX7046);
	and 	XG12545 	(WX7473,WX7474,WX7045);
	and 	XG12546 	(WX6397,WX6398,WX5783);
	and 	XG12547 	(WX6390,WX6391,WX5782);
	and 	XG12548 	(WX6383,WX6384,WX5781);
	and 	XG12549 	(WX6376,WX6377,WX5780);
	and 	XG12550 	(WX6369,WX6370,WX5779);
	and 	XG12551 	(WX6362,WX6363,WX5778);
	and 	XG12552 	(WX6355,WX6356,WX5777);
	and 	XG12553 	(WX6348,WX6349,WX5776);
	and 	XG12554 	(WX6341,WX6342,WX5775);
	and 	XG12555 	(WX6334,WX6335,WX5774);
	and 	XG12556 	(WX6327,WX6328,WX5773);
	and 	XG12557 	(WX6320,WX6321,WX5772);
	and 	XG12558 	(WX6313,WX6314,WX5771);
	and 	XG12559 	(WX6306,WX6307,WX5770);
	and 	XG12560 	(WX6299,WX6300,WX5769);
	and 	XG12561 	(WX6292,WX6293,WX5768);
	and 	XG12562 	(WX6285,WX6286,WX5767);
	and 	XG12563 	(WX6278,WX6279,WX5766);
	and 	XG12564 	(WX6271,WX6272,WX5765);
	and 	XG12565 	(WX6264,WX6265,WX5764);
	and 	XG12566 	(WX6257,WX6258,WX5763);
	and 	XG12567 	(WX6250,WX6251,WX5762);
	and 	XG12568 	(WX6243,WX6244,WX5761);
	and 	XG12569 	(WX6236,WX6237,WX5760);
	and 	XG12570 	(WX6229,WX6230,WX5759);
	and 	XG12571 	(WX6222,WX6223,WX5758);
	and 	XG12572 	(WX6215,WX6216,WX5757);
	and 	XG12573 	(WX6208,WX6209,WX5756);
	and 	XG12574 	(WX6201,WX6202,WX5755);
	and 	XG12575 	(WX6194,WX6195,WX5754);
	and 	XG12576 	(WX6187,WX6188,WX5753);
	and 	XG12577 	(WX6180,WX6181,WX5752);
	and 	XG12578 	(WX5104,WX5105,WX4490);
	and 	XG12579 	(WX5097,WX5098,WX4489);
	and 	XG12580 	(WX5090,WX5091,WX4488);
	and 	XG12581 	(WX5083,WX5084,WX4487);
	and 	XG12582 	(WX5076,WX5077,WX4486);
	and 	XG12583 	(WX5069,WX5070,WX4485);
	and 	XG12584 	(WX5062,WX5063,WX4484);
	and 	XG12585 	(WX5055,WX5056,WX4483);
	and 	XG12586 	(WX5048,WX5049,WX4482);
	and 	XG12587 	(WX5041,WX5042,WX4481);
	and 	XG12588 	(WX5034,WX5035,WX4480);
	and 	XG12589 	(WX5027,WX5028,WX4479);
	and 	XG12590 	(WX5020,WX5021,WX4478);
	and 	XG12591 	(WX5013,WX5014,WX4477);
	and 	XG12592 	(WX5006,WX5007,WX4476);
	and 	XG12593 	(WX4999,WX5000,WX4475);
	and 	XG12594 	(WX4992,WX4993,WX4474);
	and 	XG12595 	(WX4985,WX4986,WX4473);
	and 	XG12596 	(WX4978,WX4979,WX4472);
	and 	XG12597 	(WX4971,WX4972,WX4471);
	and 	XG12598 	(WX4964,WX4965,WX4470);
	and 	XG12599 	(WX4957,WX4958,WX4469);
	and 	XG12600 	(WX4950,WX4951,WX4468);
	and 	XG12601 	(WX4943,WX4944,WX4467);
	and 	XG12602 	(WX4936,WX4937,WX4466);
	and 	XG12603 	(WX4929,WX4930,WX4465);
	and 	XG12604 	(WX4922,WX4923,WX4464);
	and 	XG12605 	(WX4915,WX4916,WX4463);
	and 	XG12606 	(WX4908,WX4909,WX4462);
	and 	XG12607 	(WX4901,WX4902,WX4461);
	and 	XG12608 	(WX4894,WX4895,WX4460);
	and 	XG12609 	(WX4887,WX4888,WX4459);
	and 	XG12610 	(WX3811,WX3812,WX3197);
	and 	XG12611 	(WX3804,WX3805,WX3196);
	and 	XG12612 	(WX3797,WX3798,WX3195);
	and 	XG12613 	(WX3790,WX3791,WX3194);
	and 	XG12614 	(WX3783,WX3784,WX3193);
	and 	XG12615 	(WX3776,WX3777,WX3192);
	and 	XG12616 	(WX3769,WX3770,WX3191);
	and 	XG12617 	(WX3762,WX3763,WX3190);
	and 	XG12618 	(WX3755,WX3756,WX3189);
	and 	XG12619 	(WX3748,WX3749,WX3188);
	and 	XG12620 	(WX3741,WX3742,WX3187);
	and 	XG12621 	(WX3734,WX3735,WX3186);
	and 	XG12622 	(WX3727,WX3728,WX3185);
	and 	XG12623 	(WX3720,WX3721,WX3184);
	and 	XG12624 	(WX3713,WX3714,WX3183);
	and 	XG12625 	(WX3706,WX3707,WX3182);
	and 	XG12626 	(WX3699,WX3700,WX3181);
	and 	XG12627 	(WX3692,WX3693,WX3180);
	and 	XG12628 	(WX3685,WX3686,WX3179);
	and 	XG12629 	(WX3678,WX3679,WX3178);
	and 	XG12630 	(WX3671,WX3672,WX3177);
	and 	XG12631 	(WX3664,WX3665,WX3176);
	and 	XG12632 	(WX3657,WX3658,WX3175);
	and 	XG12633 	(WX3650,WX3651,WX3174);
	and 	XG12634 	(WX3643,WX3644,WX3173);
	and 	XG12635 	(WX3636,WX3637,WX3172);
	and 	XG12636 	(WX3629,WX3630,WX3171);
	and 	XG12637 	(WX3622,WX3623,WX3170);
	and 	XG12638 	(WX3615,WX3616,WX3169);
	and 	XG12639 	(WX3608,WX3609,WX3168);
	and 	XG12640 	(WX3601,WX3602,WX3167);
	and 	XG12641 	(WX3594,WX3595,WX3166);
	and 	XG12642 	(WX2518,WX2519,WX1904);
	and 	XG12643 	(WX2511,WX2512,WX1903);
	and 	XG12644 	(WX2504,WX2505,WX1902);
	and 	XG12645 	(WX2497,WX2498,WX1901);
	and 	XG12646 	(WX2490,WX2491,WX1900);
	and 	XG12647 	(WX2483,WX2484,WX1899);
	and 	XG12648 	(WX2476,WX2477,WX1898);
	and 	XG12649 	(WX2469,WX2470,WX1897);
	and 	XG12650 	(WX2462,WX2463,WX1896);
	and 	XG12651 	(WX2455,WX2456,WX1895);
	and 	XG12652 	(WX2448,WX2449,WX1894);
	and 	XG12653 	(WX2441,WX2442,WX1893);
	and 	XG12654 	(WX2434,WX2435,WX1892);
	and 	XG12655 	(WX2427,WX2428,WX1891);
	and 	XG12656 	(WX2420,WX2421,WX1890);
	and 	XG12657 	(WX2413,WX2414,WX1889);
	and 	XG12658 	(WX2406,WX2407,WX1888);
	and 	XG12659 	(WX2399,WX2400,WX1887);
	and 	XG12660 	(WX2392,WX2393,WX1886);
	and 	XG12661 	(WX2385,WX2386,WX1885);
	and 	XG12662 	(WX2378,WX2379,WX1884);
	and 	XG12663 	(WX2371,WX2372,WX1883);
	and 	XG12664 	(WX2364,WX2365,WX1882);
	and 	XG12665 	(WX2357,WX2358,WX1881);
	and 	XG12666 	(WX2350,WX2351,WX1880);
	and 	XG12667 	(WX2343,WX2344,WX1879);
	and 	XG12668 	(WX2336,WX2337,WX1878);
	and 	XG12669 	(WX2329,WX2330,WX1877);
	and 	XG12670 	(WX2322,WX2323,WX1876);
	and 	XG12671 	(WX2315,WX2316,WX1875);
	and 	XG12672 	(WX2308,WX2309,WX1874);
	and 	XG12673 	(WX2301,WX2302,WX1873);
	and 	XG12674 	(WX1225,WX1226,WX611);
	and 	XG12675 	(WX1218,WX1219,WX610);
	and 	XG12676 	(WX1211,WX1212,WX609);
	and 	XG12677 	(WX1204,WX1205,WX608);
	and 	XG12678 	(WX1197,WX1198,WX607);
	and 	XG12679 	(WX1190,WX1191,WX606);
	and 	XG12680 	(WX1183,WX1184,WX605);
	and 	XG12681 	(WX1176,WX1177,WX604);
	and 	XG12682 	(WX1169,WX1170,WX603);
	and 	XG12683 	(WX1162,WX1163,WX602);
	and 	XG12684 	(WX1155,WX1156,WX601);
	and 	XG12685 	(WX1148,WX1149,WX600);
	and 	XG12686 	(WX1141,WX1142,WX599);
	and 	XG12687 	(WX1134,WX1135,WX598);
	and 	XG12688 	(WX1127,WX1128,WX597);
	and 	XG12689 	(WX1120,WX1121,WX596);
	and 	XG12690 	(WX1113,WX1114,WX595);
	and 	XG12691 	(WX1106,WX1107,WX594);
	and 	XG12692 	(WX1099,WX1100,WX593);
	and 	XG12693 	(WX1092,WX1093,WX592);
	and 	XG12694 	(WX1085,WX1086,WX591);
	and 	XG12695 	(WX1078,WX1079,WX590);
	and 	XG12696 	(WX1071,WX1072,WX589);
	and 	XG12697 	(WX1064,WX1065,WX588);
	and 	XG12698 	(WX1057,WX1058,WX587);
	and 	XG12699 	(WX1050,WX1051,WX586);
	and 	XG12700 	(WX1043,WX1044,WX585);
	and 	XG12701 	(WX1036,WX1037,WX584);
	and 	XG12702 	(WX1029,WX1030,WX583);
	and 	XG12703 	(WX1022,WX1023,WX582);
	and 	XG12704 	(WX1015,WX1016,WX581);
	and 	XG12705 	(WX1008,WX1009,WX580);
	nand 	XG12706 	(II3052,WX485,WX580);
	nand 	XG12707 	(II3065,WX487,WX581);
	nand 	XG12708 	(II3078,WX489,WX582);
	nand 	XG12709 	(II3091,WX491,WX583);
	nand 	XG12710 	(II3104,WX493,WX584);
	nand 	XG12711 	(II3117,WX495,WX585);
	nand 	XG12712 	(II3130,WX497,WX586);
	nand 	XG12713 	(II3143,WX499,WX587);
	nand 	XG12714 	(II3156,WX501,WX588);
	nand 	XG12715 	(II3169,WX503,WX589);
	nand 	XG12716 	(II3182,WX505,WX590);
	nand 	XG12717 	(II3195,WX507,WX591);
	nand 	XG12718 	(II3208,WX509,WX592);
	nand 	XG12719 	(II3221,WX511,WX593);
	nand 	XG12720 	(II3234,WX513,WX594);
	nand 	XG12721 	(II3247,WX515,WX595);
	nand 	XG12722 	(II3260,WX517,WX596);
	nand 	XG12723 	(II3273,WX519,WX597);
	nand 	XG12724 	(II3286,WX521,WX598);
	nand 	XG12725 	(II3299,WX523,WX599);
	nand 	XG12726 	(II3312,WX525,WX600);
	nand 	XG12727 	(II3325,WX527,WX601);
	nand 	XG12728 	(II3338,WX529,WX602);
	nand 	XG12729 	(II3351,WX531,WX603);
	nand 	XG12730 	(II3364,WX533,WX604);
	nand 	XG12731 	(II3377,WX535,WX605);
	nand 	XG12732 	(II3390,WX537,WX606);
	nand 	XG12733 	(II3403,WX539,WX607);
	nand 	XG12734 	(II3416,WX541,WX608);
	nand 	XG12735 	(II3429,WX543,WX609);
	nand 	XG12736 	(II3442,WX545,WX610);
	nand 	XG12737 	(II3455,WX547,WX611);
	nand 	XG12738 	(II7057,WX1778,WX1873);
	nand 	XG12739 	(II7070,WX1780,WX1874);
	nand 	XG12740 	(II7083,WX1782,WX1875);
	nand 	XG12741 	(II7096,WX1784,WX1876);
	nand 	XG12742 	(II7109,WX1786,WX1877);
	nand 	XG12743 	(II7122,WX1788,WX1878);
	nand 	XG12744 	(II7135,WX1790,WX1879);
	nand 	XG12745 	(II7148,WX1792,WX1880);
	nand 	XG12746 	(II7161,WX1794,WX1881);
	nand 	XG12747 	(II7174,WX1796,WX1882);
	nand 	XG12748 	(II7187,WX1798,WX1883);
	nand 	XG12749 	(II7200,WX1800,WX1884);
	nand 	XG12750 	(II7213,WX1802,WX1885);
	nand 	XG12751 	(II7226,WX1804,WX1886);
	nand 	XG12752 	(II7239,WX1806,WX1887);
	nand 	XG12753 	(II7252,WX1808,WX1888);
	nand 	XG12754 	(II7265,WX1810,WX1889);
	nand 	XG12755 	(II7278,WX1812,WX1890);
	nand 	XG12756 	(II7291,WX1814,WX1891);
	nand 	XG12757 	(II7304,WX1816,WX1892);
	nand 	XG12758 	(II7317,WX1818,WX1893);
	nand 	XG12759 	(II7330,WX1820,WX1894);
	nand 	XG12760 	(II7343,WX1822,WX1895);
	nand 	XG12761 	(II7356,WX1824,WX1896);
	nand 	XG12762 	(II7369,WX1826,WX1897);
	nand 	XG12763 	(II7382,WX1828,WX1898);
	nand 	XG12764 	(II7395,WX1830,WX1899);
	nand 	XG12765 	(II7408,WX1832,WX1900);
	nand 	XG12766 	(II7421,WX1834,WX1901);
	nand 	XG12767 	(II7434,WX1836,WX1902);
	nand 	XG12768 	(II7447,WX1838,WX1903);
	nand 	XG12769 	(II7460,WX1840,WX1904);
	nand 	XG12770 	(II11062,WX3071,WX3166);
	nand 	XG12771 	(II11075,WX3073,WX3167);
	nand 	XG12772 	(II11088,WX3075,WX3168);
	nand 	XG12773 	(II11101,WX3077,WX3169);
	nand 	XG12774 	(II11114,WX3079,WX3170);
	nand 	XG12775 	(II11127,WX3081,WX3171);
	nand 	XG12776 	(II11140,WX3083,WX3172);
	nand 	XG12777 	(II11153,WX3085,WX3173);
	nand 	XG12778 	(II11166,WX3087,WX3174);
	nand 	XG12779 	(II11179,WX3089,WX3175);
	nand 	XG12780 	(II11192,WX3091,WX3176);
	nand 	XG12781 	(II11205,WX3093,WX3177);
	nand 	XG12782 	(II11218,WX3095,WX3178);
	nand 	XG12783 	(II11231,WX3097,WX3179);
	nand 	XG12784 	(II11244,WX3099,WX3180);
	nand 	XG12785 	(II11257,WX3101,WX3181);
	nand 	XG12786 	(II11270,WX3103,WX3182);
	nand 	XG12787 	(II11283,WX3105,WX3183);
	nand 	XG12788 	(II11296,WX3107,WX3184);
	nand 	XG12789 	(II11309,WX3109,WX3185);
	nand 	XG12790 	(II11322,WX3111,WX3186);
	nand 	XG12791 	(II11335,WX3113,WX3187);
	nand 	XG12792 	(II11348,WX3115,WX3188);
	nand 	XG12793 	(II11361,WX3117,WX3189);
	nand 	XG12794 	(II11374,WX3119,WX3190);
	nand 	XG12795 	(II11387,WX3121,WX3191);
	nand 	XG12796 	(II11400,WX3123,WX3192);
	nand 	XG12797 	(II11413,WX3125,WX3193);
	nand 	XG12798 	(II11426,WX3127,WX3194);
	nand 	XG12799 	(II11439,WX3129,WX3195);
	nand 	XG12800 	(II11452,WX3131,WX3196);
	nand 	XG12801 	(II11465,WX3133,WX3197);
	nand 	XG12802 	(II15067,WX4364,WX4459);
	nand 	XG12803 	(II15080,WX4366,WX4460);
	nand 	XG12804 	(II15093,WX4368,WX4461);
	nand 	XG12805 	(II15106,WX4370,WX4462);
	nand 	XG12806 	(II15119,WX4372,WX4463);
	nand 	XG12807 	(II15132,WX4374,WX4464);
	nand 	XG12808 	(II15145,WX4376,WX4465);
	nand 	XG12809 	(II15158,WX4378,WX4466);
	nand 	XG12810 	(II15171,WX4380,WX4467);
	nand 	XG12811 	(II15184,WX4382,WX4468);
	nand 	XG12812 	(II15197,WX4384,WX4469);
	nand 	XG12813 	(II15210,WX4386,WX4470);
	nand 	XG12814 	(II15223,WX4388,WX4471);
	nand 	XG12815 	(II15236,WX4390,WX4472);
	nand 	XG12816 	(II15249,WX4392,WX4473);
	nand 	XG12817 	(II15262,WX4394,WX4474);
	nand 	XG12818 	(II15275,WX4396,WX4475);
	nand 	XG12819 	(II15288,WX4398,WX4476);
	nand 	XG12820 	(II15301,WX4400,WX4477);
	nand 	XG12821 	(II15314,WX4402,WX4478);
	nand 	XG12822 	(II15327,WX4404,WX4479);
	nand 	XG12823 	(II15340,WX4406,WX4480);
	nand 	XG12824 	(II15353,WX4408,WX4481);
	nand 	XG12825 	(II15366,WX4410,WX4482);
	nand 	XG12826 	(II15379,WX4412,WX4483);
	nand 	XG12827 	(II15392,WX4414,WX4484);
	nand 	XG12828 	(II15405,WX4416,WX4485);
	nand 	XG12829 	(II15418,WX4418,WX4486);
	nand 	XG12830 	(II15431,WX4420,WX4487);
	nand 	XG12831 	(II15444,WX4422,WX4488);
	nand 	XG12832 	(II15457,WX4424,WX4489);
	nand 	XG12833 	(II15470,WX4426,WX4490);
	nand 	XG12834 	(II19072,WX5657,WX5752);
	nand 	XG12835 	(II19085,WX5659,WX5753);
	nand 	XG12836 	(II19098,WX5661,WX5754);
	nand 	XG12837 	(II19111,WX5663,WX5755);
	nand 	XG12838 	(II19124,WX5665,WX5756);
	nand 	XG12839 	(II19137,WX5667,WX5757);
	nand 	XG12840 	(II19150,WX5669,WX5758);
	nand 	XG12841 	(II19163,WX5671,WX5759);
	nand 	XG12842 	(II19176,WX5673,WX5760);
	nand 	XG12843 	(II19189,WX5675,WX5761);
	nand 	XG12844 	(II19202,WX5677,WX5762);
	nand 	XG12845 	(II19215,WX5679,WX5763);
	nand 	XG12846 	(II19228,WX5681,WX5764);
	nand 	XG12847 	(II19241,WX5683,WX5765);
	nand 	XG12848 	(II19254,WX5685,WX5766);
	nand 	XG12849 	(II19267,WX5687,WX5767);
	nand 	XG12850 	(II19280,WX5689,WX5768);
	nand 	XG12851 	(II19293,WX5691,WX5769);
	nand 	XG12852 	(II19306,WX5693,WX5770);
	nand 	XG12853 	(II19319,WX5695,WX5771);
	nand 	XG12854 	(II19332,WX5697,WX5772);
	nand 	XG12855 	(II19345,WX5699,WX5773);
	nand 	XG12856 	(II19358,WX5701,WX5774);
	nand 	XG12857 	(II19371,WX5703,WX5775);
	nand 	XG12858 	(II19384,WX5705,WX5776);
	nand 	XG12859 	(II19397,WX5707,WX5777);
	nand 	XG12860 	(II19410,WX5709,WX5778);
	nand 	XG12861 	(II19423,WX5711,WX5779);
	nand 	XG12862 	(II19436,WX5713,WX5780);
	nand 	XG12863 	(II19449,WX5715,WX5781);
	nand 	XG12864 	(II19462,WX5717,WX5782);
	nand 	XG12865 	(II19475,WX5719,WX5783);
	nand 	XG12866 	(II23077,WX6950,WX7045);
	nand 	XG12867 	(II23090,WX6952,WX7046);
	nand 	XG12868 	(II23103,WX6954,WX7047);
	nand 	XG12869 	(II23116,WX6956,WX7048);
	nand 	XG12870 	(II23129,WX6958,WX7049);
	nand 	XG12871 	(II23142,WX6960,WX7050);
	nand 	XG12872 	(II23155,WX6962,WX7051);
	nand 	XG12873 	(II23168,WX6964,WX7052);
	nand 	XG12874 	(II23181,WX6966,WX7053);
	nand 	XG12875 	(II23194,WX6968,WX7054);
	nand 	XG12876 	(II23207,WX6970,WX7055);
	nand 	XG12877 	(II23220,WX6972,WX7056);
	nand 	XG12878 	(II23233,WX6974,WX7057);
	nand 	XG12879 	(II23246,WX6976,WX7058);
	nand 	XG12880 	(II23259,WX6978,WX7059);
	nand 	XG12881 	(II23272,WX6980,WX7060);
	nand 	XG12882 	(II23285,WX6982,WX7061);
	nand 	XG12883 	(II23298,WX6984,WX7062);
	nand 	XG12884 	(II23311,WX6986,WX7063);
	nand 	XG12885 	(II23324,WX6988,WX7064);
	nand 	XG12886 	(II23337,WX6990,WX7065);
	nand 	XG12887 	(II23350,WX6992,WX7066);
	nand 	XG12888 	(II23363,WX6994,WX7067);
	nand 	XG12889 	(II23376,WX6996,WX7068);
	nand 	XG12890 	(II23389,WX6998,WX7069);
	nand 	XG12891 	(II23402,WX7000,WX7070);
	nand 	XG12892 	(II23415,WX7002,WX7071);
	nand 	XG12893 	(II23428,WX7004,WX7072);
	nand 	XG12894 	(II23441,WX7006,WX7073);
	nand 	XG12895 	(II23454,WX7008,WX7074);
	nand 	XG12896 	(II23467,WX7010,WX7075);
	nand 	XG12897 	(II23480,WX7012,WX7076);
	nand 	XG12898 	(II27082,WX8243,WX8338);
	nand 	XG12899 	(II27095,WX8245,WX8339);
	nand 	XG12900 	(II27108,WX8247,WX8340);
	nand 	XG12901 	(II27121,WX8249,WX8341);
	nand 	XG12902 	(II27134,WX8251,WX8342);
	nand 	XG12903 	(II27147,WX8253,WX8343);
	nand 	XG12904 	(II27160,WX8255,WX8344);
	nand 	XG12905 	(II27173,WX8257,WX8345);
	nand 	XG12906 	(II27186,WX8259,WX8346);
	nand 	XG12907 	(II27199,WX8261,WX8347);
	nand 	XG12908 	(II27212,WX8263,WX8348);
	nand 	XG12909 	(II27225,WX8265,WX8349);
	nand 	XG12910 	(II27238,WX8267,WX8350);
	nand 	XG12911 	(II27251,WX8269,WX8351);
	nand 	XG12912 	(II27264,WX8271,WX8352);
	nand 	XG12913 	(II27277,WX8273,WX8353);
	nand 	XG12914 	(II27290,WX8275,WX8354);
	nand 	XG12915 	(II27303,WX8277,WX8355);
	nand 	XG12916 	(II27316,WX8279,WX8356);
	nand 	XG12917 	(II27329,WX8281,WX8357);
	nand 	XG12918 	(II27342,WX8283,WX8358);
	nand 	XG12919 	(II27355,WX8285,WX8359);
	nand 	XG12920 	(II27368,WX8287,WX8360);
	nand 	XG12921 	(II27381,WX8289,WX8361);
	nand 	XG12922 	(II27394,WX8291,WX8362);
	nand 	XG12923 	(II27407,WX8293,WX8363);
	nand 	XG12924 	(II27420,WX8295,WX8364);
	nand 	XG12925 	(II27433,WX8297,WX8365);
	nand 	XG12926 	(II27446,WX8299,WX8366);
	nand 	XG12927 	(II27459,WX8301,WX8367);
	nand 	XG12928 	(II27472,WX8303,WX8368);
	nand 	XG12929 	(II27485,WX8305,WX8369);
	nand 	XG12930 	(II31087,WX9536,WX9631);
	nand 	XG12931 	(II31100,WX9538,WX9632);
	nand 	XG12932 	(II31113,WX9540,WX9633);
	nand 	XG12933 	(II31126,WX9542,WX9634);
	nand 	XG12934 	(II31139,WX9544,WX9635);
	nand 	XG12935 	(II31152,WX9546,WX9636);
	nand 	XG12936 	(II31165,WX9548,WX9637);
	nand 	XG12937 	(II31178,WX9550,WX9638);
	nand 	XG12938 	(II31191,WX9552,WX9639);
	nand 	XG12939 	(II31204,WX9554,WX9640);
	nand 	XG12940 	(II31217,WX9556,WX9641);
	nand 	XG12941 	(II31230,WX9558,WX9642);
	nand 	XG12942 	(II31243,WX9560,WX9643);
	nand 	XG12943 	(II31256,WX9562,WX9644);
	nand 	XG12944 	(II31269,WX9564,WX9645);
	nand 	XG12945 	(II31282,WX9566,WX9646);
	nand 	XG12946 	(II31295,WX9568,WX9647);
	nand 	XG12947 	(II31308,WX9570,WX9648);
	nand 	XG12948 	(II31321,WX9572,WX9649);
	nand 	XG12949 	(II31334,WX9574,WX9650);
	nand 	XG12950 	(II31347,WX9576,WX9651);
	nand 	XG12951 	(II31360,WX9578,WX9652);
	nand 	XG12952 	(II31373,WX9580,WX9653);
	nand 	XG12953 	(II31386,WX9582,WX9654);
	nand 	XG12954 	(II31399,WX9584,WX9655);
	nand 	XG12955 	(II31412,WX9586,WX9656);
	nand 	XG12956 	(II31425,WX9588,WX9657);
	nand 	XG12957 	(II31438,WX9590,WX9658);
	nand 	XG12958 	(II31451,WX9592,WX9659);
	nand 	XG12959 	(II31464,WX9594,WX9660);
	nand 	XG12960 	(II31477,WX9596,WX9661);
	nand 	XG12961 	(II31490,WX9598,WX9662);
	nand 	XG12962 	(II35092,WX10829,WX10924);
	nand 	XG12963 	(II35105,WX10831,WX10925);
	nand 	XG12964 	(II35118,WX10833,WX10926);
	nand 	XG12965 	(II35131,WX10835,WX10927);
	nand 	XG12966 	(II35144,WX10837,WX10928);
	nand 	XG12967 	(II35157,WX10839,WX10929);
	nand 	XG12968 	(II35170,WX10841,WX10930);
	nand 	XG12969 	(II35183,WX10843,WX10931);
	nand 	XG12970 	(II35196,WX10845,WX10932);
	nand 	XG12971 	(II35209,WX10847,WX10933);
	nand 	XG12972 	(II35222,WX10849,WX10934);
	nand 	XG12973 	(II35235,WX10851,WX10935);
	nand 	XG12974 	(II35248,WX10853,WX10936);
	nand 	XG12975 	(II35261,WX10855,WX10937);
	nand 	XG12976 	(II35274,WX10857,WX10938);
	nand 	XG12977 	(II35287,WX10859,WX10939);
	nand 	XG12978 	(II35300,WX10861,WX10940);
	nand 	XG12979 	(II35313,WX10863,WX10941);
	nand 	XG12980 	(II35326,WX10865,WX10942);
	nand 	XG12981 	(II35339,WX10867,WX10943);
	nand 	XG12982 	(II35352,WX10869,WX10944);
	nand 	XG12983 	(II35365,WX10871,WX10945);
	nand 	XG12984 	(II35378,WX10873,WX10946);
	nand 	XG12985 	(II35391,WX10875,WX10947);
	nand 	XG12986 	(II35404,WX10877,WX10948);
	nand 	XG12987 	(II35417,WX10879,WX10949);
	nand 	XG12988 	(II35430,WX10881,WX10950);
	nand 	XG12989 	(II35443,WX10883,WX10951);
	nand 	XG12990 	(II35456,WX10885,WX10952);
	nand 	XG12991 	(II35469,WX10887,WX10953);
	nand 	XG12992 	(II35482,WX10889,WX10954);
	nand 	XG12993 	(II35495,WX10891,WX10955);
	nand 	XG12994 	(II35496,II35495,WX10955);
	nand 	XG12995 	(II35483,II35482,WX10954);
	nand 	XG12996 	(II35470,II35469,WX10953);
	nand 	XG12997 	(II35457,II35456,WX10952);
	nand 	XG12998 	(II35444,II35443,WX10951);
	nand 	XG12999 	(II35431,II35430,WX10950);
	nand 	XG13000 	(II35418,II35417,WX10949);
	nand 	XG13001 	(II35405,II35404,WX10948);
	nand 	XG13002 	(II35392,II35391,WX10947);
	nand 	XG13003 	(II35379,II35378,WX10946);
	nand 	XG13004 	(II35366,II35365,WX10945);
	nand 	XG13005 	(II35353,II35352,WX10944);
	nand 	XG13006 	(II35340,II35339,WX10943);
	nand 	XG13007 	(II35327,II35326,WX10942);
	nand 	XG13008 	(II35314,II35313,WX10941);
	nand 	XG13009 	(II35301,II35300,WX10940);
	nand 	XG13010 	(II35288,II35287,WX10939);
	nand 	XG13011 	(II35275,II35274,WX10938);
	nand 	XG13012 	(II35262,II35261,WX10937);
	nand 	XG13013 	(II35249,II35248,WX10936);
	nand 	XG13014 	(II35236,II35235,WX10935);
	nand 	XG13015 	(II35223,II35222,WX10934);
	nand 	XG13016 	(II35210,II35209,WX10933);
	nand 	XG13017 	(II35197,II35196,WX10932);
	nand 	XG13018 	(II35184,II35183,WX10931);
	nand 	XG13019 	(II35171,II35170,WX10930);
	nand 	XG13020 	(II35158,II35157,WX10929);
	nand 	XG13021 	(II35145,II35144,WX10928);
	nand 	XG13022 	(II35132,II35131,WX10927);
	nand 	XG13023 	(II35119,II35118,WX10926);
	nand 	XG13024 	(II35106,II35105,WX10925);
	nand 	XG13025 	(II35093,II35092,WX10924);
	nand 	XG13026 	(II31491,II31490,WX9662);
	nand 	XG13027 	(II31478,II31477,WX9661);
	nand 	XG13028 	(II31465,II31464,WX9660);
	nand 	XG13029 	(II31452,II31451,WX9659);
	nand 	XG13030 	(II31439,II31438,WX9658);
	nand 	XG13031 	(II31426,II31425,WX9657);
	nand 	XG13032 	(II31413,II31412,WX9656);
	nand 	XG13033 	(II31400,II31399,WX9655);
	nand 	XG13034 	(II31387,II31386,WX9654);
	nand 	XG13035 	(II31374,II31373,WX9653);
	nand 	XG13036 	(II31361,II31360,WX9652);
	nand 	XG13037 	(II31348,II31347,WX9651);
	nand 	XG13038 	(II31335,II31334,WX9650);
	nand 	XG13039 	(II31322,II31321,WX9649);
	nand 	XG13040 	(II31309,II31308,WX9648);
	nand 	XG13041 	(II31296,II31295,WX9647);
	nand 	XG13042 	(II31283,II31282,WX9646);
	nand 	XG13043 	(II31270,II31269,WX9645);
	nand 	XG13044 	(II31257,II31256,WX9644);
	nand 	XG13045 	(II31244,II31243,WX9643);
	nand 	XG13046 	(II31231,II31230,WX9642);
	nand 	XG13047 	(II31218,II31217,WX9641);
	nand 	XG13048 	(II31205,II31204,WX9640);
	nand 	XG13049 	(II31192,II31191,WX9639);
	nand 	XG13050 	(II31179,II31178,WX9638);
	nand 	XG13051 	(II31166,II31165,WX9637);
	nand 	XG13052 	(II31153,II31152,WX9636);
	nand 	XG13053 	(II31140,II31139,WX9635);
	nand 	XG13054 	(II31127,II31126,WX9634);
	nand 	XG13055 	(II31114,II31113,WX9633);
	nand 	XG13056 	(II31101,II31100,WX9632);
	nand 	XG13057 	(II31088,II31087,WX9631);
	nand 	XG13058 	(II27486,II27485,WX8369);
	nand 	XG13059 	(II27473,II27472,WX8368);
	nand 	XG13060 	(II27460,II27459,WX8367);
	nand 	XG13061 	(II27447,II27446,WX8366);
	nand 	XG13062 	(II27434,II27433,WX8365);
	nand 	XG13063 	(II27421,II27420,WX8364);
	nand 	XG13064 	(II27408,II27407,WX8363);
	nand 	XG13065 	(II27395,II27394,WX8362);
	nand 	XG13066 	(II27382,II27381,WX8361);
	nand 	XG13067 	(II27369,II27368,WX8360);
	nand 	XG13068 	(II27356,II27355,WX8359);
	nand 	XG13069 	(II27343,II27342,WX8358);
	nand 	XG13070 	(II27330,II27329,WX8357);
	nand 	XG13071 	(II27317,II27316,WX8356);
	nand 	XG13072 	(II27304,II27303,WX8355);
	nand 	XG13073 	(II27291,II27290,WX8354);
	nand 	XG13074 	(II27278,II27277,WX8353);
	nand 	XG13075 	(II27265,II27264,WX8352);
	nand 	XG13076 	(II27252,II27251,WX8351);
	nand 	XG13077 	(II27239,II27238,WX8350);
	nand 	XG13078 	(II27226,II27225,WX8349);
	nand 	XG13079 	(II27213,II27212,WX8348);
	nand 	XG13080 	(II27200,II27199,WX8347);
	nand 	XG13081 	(II27187,II27186,WX8346);
	nand 	XG13082 	(II27174,II27173,WX8345);
	nand 	XG13083 	(II27161,II27160,WX8344);
	nand 	XG13084 	(II27148,II27147,WX8343);
	nand 	XG13085 	(II27135,II27134,WX8342);
	nand 	XG13086 	(II27122,II27121,WX8341);
	nand 	XG13087 	(II27109,II27108,WX8340);
	nand 	XG13088 	(II27096,II27095,WX8339);
	nand 	XG13089 	(II27083,II27082,WX8338);
	nand 	XG13090 	(II23481,II23480,WX7076);
	nand 	XG13091 	(II23468,II23467,WX7075);
	nand 	XG13092 	(II23455,II23454,WX7074);
	nand 	XG13093 	(II23442,II23441,WX7073);
	nand 	XG13094 	(II23429,II23428,WX7072);
	nand 	XG13095 	(II23416,II23415,WX7071);
	nand 	XG13096 	(II23403,II23402,WX7070);
	nand 	XG13097 	(II23390,II23389,WX7069);
	nand 	XG13098 	(II23377,II23376,WX7068);
	nand 	XG13099 	(II23364,II23363,WX7067);
	nand 	XG13100 	(II23351,II23350,WX7066);
	nand 	XG13101 	(II23338,II23337,WX7065);
	nand 	XG13102 	(II23325,II23324,WX7064);
	nand 	XG13103 	(II23312,II23311,WX7063);
	nand 	XG13104 	(II23299,II23298,WX7062);
	nand 	XG13105 	(II23286,II23285,WX7061);
	nand 	XG13106 	(II23273,II23272,WX7060);
	nand 	XG13107 	(II23260,II23259,WX7059);
	nand 	XG13108 	(II23247,II23246,WX7058);
	nand 	XG13109 	(II23234,II23233,WX7057);
	nand 	XG13110 	(II23221,II23220,WX7056);
	nand 	XG13111 	(II23208,II23207,WX7055);
	nand 	XG13112 	(II23195,II23194,WX7054);
	nand 	XG13113 	(II23182,II23181,WX7053);
	nand 	XG13114 	(II23169,II23168,WX7052);
	nand 	XG13115 	(II23156,II23155,WX7051);
	nand 	XG13116 	(II23143,II23142,WX7050);
	nand 	XG13117 	(II23130,II23129,WX7049);
	nand 	XG13118 	(II23117,II23116,WX7048);
	nand 	XG13119 	(II23104,II23103,WX7047);
	nand 	XG13120 	(II23091,II23090,WX7046);
	nand 	XG13121 	(II23078,II23077,WX7045);
	nand 	XG13122 	(II19476,II19475,WX5783);
	nand 	XG13123 	(II19463,II19462,WX5782);
	nand 	XG13124 	(II19450,II19449,WX5781);
	nand 	XG13125 	(II19437,II19436,WX5780);
	nand 	XG13126 	(II19424,II19423,WX5779);
	nand 	XG13127 	(II19411,II19410,WX5778);
	nand 	XG13128 	(II19398,II19397,WX5777);
	nand 	XG13129 	(II19385,II19384,WX5776);
	nand 	XG13130 	(II19372,II19371,WX5775);
	nand 	XG13131 	(II19359,II19358,WX5774);
	nand 	XG13132 	(II19346,II19345,WX5773);
	nand 	XG13133 	(II19333,II19332,WX5772);
	nand 	XG13134 	(II19320,II19319,WX5771);
	nand 	XG13135 	(II19307,II19306,WX5770);
	nand 	XG13136 	(II19294,II19293,WX5769);
	nand 	XG13137 	(II19281,II19280,WX5768);
	nand 	XG13138 	(II19268,II19267,WX5767);
	nand 	XG13139 	(II19255,II19254,WX5766);
	nand 	XG13140 	(II19242,II19241,WX5765);
	nand 	XG13141 	(II19229,II19228,WX5764);
	nand 	XG13142 	(II19216,II19215,WX5763);
	nand 	XG13143 	(II19203,II19202,WX5762);
	nand 	XG13144 	(II19190,II19189,WX5761);
	nand 	XG13145 	(II19177,II19176,WX5760);
	nand 	XG13146 	(II19164,II19163,WX5759);
	nand 	XG13147 	(II19151,II19150,WX5758);
	nand 	XG13148 	(II19138,II19137,WX5757);
	nand 	XG13149 	(II19125,II19124,WX5756);
	nand 	XG13150 	(II19112,II19111,WX5755);
	nand 	XG13151 	(II19099,II19098,WX5754);
	nand 	XG13152 	(II19086,II19085,WX5753);
	nand 	XG13153 	(II19073,II19072,WX5752);
	nand 	XG13154 	(II15471,II15470,WX4490);
	nand 	XG13155 	(II15458,II15457,WX4489);
	nand 	XG13156 	(II15445,II15444,WX4488);
	nand 	XG13157 	(II15432,II15431,WX4487);
	nand 	XG13158 	(II15419,II15418,WX4486);
	nand 	XG13159 	(II15406,II15405,WX4485);
	nand 	XG13160 	(II15393,II15392,WX4484);
	nand 	XG13161 	(II15380,II15379,WX4483);
	nand 	XG13162 	(II15367,II15366,WX4482);
	nand 	XG13163 	(II15354,II15353,WX4481);
	nand 	XG13164 	(II15341,II15340,WX4480);
	nand 	XG13165 	(II15328,II15327,WX4479);
	nand 	XG13166 	(II15315,II15314,WX4478);
	nand 	XG13167 	(II15302,II15301,WX4477);
	nand 	XG13168 	(II15289,II15288,WX4476);
	nand 	XG13169 	(II15276,II15275,WX4475);
	nand 	XG13170 	(II15263,II15262,WX4474);
	nand 	XG13171 	(II15250,II15249,WX4473);
	nand 	XG13172 	(II15237,II15236,WX4472);
	nand 	XG13173 	(II15224,II15223,WX4471);
	nand 	XG13174 	(II15211,II15210,WX4470);
	nand 	XG13175 	(II15198,II15197,WX4469);
	nand 	XG13176 	(II15185,II15184,WX4468);
	nand 	XG13177 	(II15172,II15171,WX4467);
	nand 	XG13178 	(II15159,II15158,WX4466);
	nand 	XG13179 	(II15146,II15145,WX4465);
	nand 	XG13180 	(II15133,II15132,WX4464);
	nand 	XG13181 	(II15120,II15119,WX4463);
	nand 	XG13182 	(II15107,II15106,WX4462);
	nand 	XG13183 	(II15094,II15093,WX4461);
	nand 	XG13184 	(II15081,II15080,WX4460);
	nand 	XG13185 	(II15068,II15067,WX4459);
	nand 	XG13186 	(II11466,II11465,WX3197);
	nand 	XG13187 	(II11453,II11452,WX3196);
	nand 	XG13188 	(II11440,II11439,WX3195);
	nand 	XG13189 	(II11427,II11426,WX3194);
	nand 	XG13190 	(II11414,II11413,WX3193);
	nand 	XG13191 	(II11401,II11400,WX3192);
	nand 	XG13192 	(II11388,II11387,WX3191);
	nand 	XG13193 	(II11375,II11374,WX3190);
	nand 	XG13194 	(II11362,II11361,WX3189);
	nand 	XG13195 	(II11349,II11348,WX3188);
	nand 	XG13196 	(II11336,II11335,WX3187);
	nand 	XG13197 	(II11323,II11322,WX3186);
	nand 	XG13198 	(II11310,II11309,WX3185);
	nand 	XG13199 	(II11297,II11296,WX3184);
	nand 	XG13200 	(II11284,II11283,WX3183);
	nand 	XG13201 	(II11271,II11270,WX3182);
	nand 	XG13202 	(II11258,II11257,WX3181);
	nand 	XG13203 	(II11245,II11244,WX3180);
	nand 	XG13204 	(II11232,II11231,WX3179);
	nand 	XG13205 	(II11219,II11218,WX3178);
	nand 	XG13206 	(II11206,II11205,WX3177);
	nand 	XG13207 	(II11193,II11192,WX3176);
	nand 	XG13208 	(II11180,II11179,WX3175);
	nand 	XG13209 	(II11167,II11166,WX3174);
	nand 	XG13210 	(II11154,II11153,WX3173);
	nand 	XG13211 	(II11141,II11140,WX3172);
	nand 	XG13212 	(II11128,II11127,WX3171);
	nand 	XG13213 	(II11115,II11114,WX3170);
	nand 	XG13214 	(II11102,II11101,WX3169);
	nand 	XG13215 	(II11089,II11088,WX3168);
	nand 	XG13216 	(II11076,II11075,WX3167);
	nand 	XG13217 	(II11063,II11062,WX3166);
	nand 	XG13218 	(II7461,II7460,WX1904);
	nand 	XG13219 	(II7448,II7447,WX1903);
	nand 	XG13220 	(II7435,II7434,WX1902);
	nand 	XG13221 	(II7422,II7421,WX1901);
	nand 	XG13222 	(II7409,II7408,WX1900);
	nand 	XG13223 	(II7396,II7395,WX1899);
	nand 	XG13224 	(II7383,II7382,WX1898);
	nand 	XG13225 	(II7370,II7369,WX1897);
	nand 	XG13226 	(II7357,II7356,WX1896);
	nand 	XG13227 	(II7344,II7343,WX1895);
	nand 	XG13228 	(II7331,II7330,WX1894);
	nand 	XG13229 	(II7318,II7317,WX1893);
	nand 	XG13230 	(II7305,II7304,WX1892);
	nand 	XG13231 	(II7292,II7291,WX1891);
	nand 	XG13232 	(II7279,II7278,WX1890);
	nand 	XG13233 	(II7266,II7265,WX1889);
	nand 	XG13234 	(II7253,II7252,WX1888);
	nand 	XG13235 	(II7240,II7239,WX1887);
	nand 	XG13236 	(II7227,II7226,WX1886);
	nand 	XG13237 	(II7214,II7213,WX1885);
	nand 	XG13238 	(II7201,II7200,WX1884);
	nand 	XG13239 	(II7188,II7187,WX1883);
	nand 	XG13240 	(II7175,II7174,WX1882);
	nand 	XG13241 	(II7162,II7161,WX1881);
	nand 	XG13242 	(II7149,II7148,WX1880);
	nand 	XG13243 	(II7136,II7135,WX1879);
	nand 	XG13244 	(II7123,II7122,WX1878);
	nand 	XG13245 	(II7110,II7109,WX1877);
	nand 	XG13246 	(II7097,II7096,WX1876);
	nand 	XG13247 	(II7084,II7083,WX1875);
	nand 	XG13248 	(II7071,II7070,WX1874);
	nand 	XG13249 	(II7058,II7057,WX1873);
	nand 	XG13250 	(II3456,II3455,WX611);
	nand 	XG13251 	(II3443,II3442,WX610);
	nand 	XG13252 	(II3430,II3429,WX609);
	nand 	XG13253 	(II3417,II3416,WX608);
	nand 	XG13254 	(II3404,II3403,WX607);
	nand 	XG13255 	(II3391,II3390,WX606);
	nand 	XG13256 	(II3378,II3377,WX605);
	nand 	XG13257 	(II3365,II3364,WX604);
	nand 	XG13258 	(II3352,II3351,WX603);
	nand 	XG13259 	(II3339,II3338,WX602);
	nand 	XG13260 	(II3326,II3325,WX601);
	nand 	XG13261 	(II3313,II3312,WX600);
	nand 	XG13262 	(II3300,II3299,WX599);
	nand 	XG13263 	(II3287,II3286,WX598);
	nand 	XG13264 	(II3274,II3273,WX597);
	nand 	XG13265 	(II3261,II3260,WX596);
	nand 	XG13266 	(II3248,II3247,WX595);
	nand 	XG13267 	(II3235,II3234,WX594);
	nand 	XG13268 	(II3222,II3221,WX593);
	nand 	XG13269 	(II3209,II3208,WX592);
	nand 	XG13270 	(II3196,II3195,WX591);
	nand 	XG13271 	(II3183,II3182,WX590);
	nand 	XG13272 	(II3170,II3169,WX589);
	nand 	XG13273 	(II3157,II3156,WX588);
	nand 	XG13274 	(II3144,II3143,WX587);
	nand 	XG13275 	(II3131,II3130,WX586);
	nand 	XG13276 	(II3118,II3117,WX585);
	nand 	XG13277 	(II3105,II3104,WX584);
	nand 	XG13278 	(II3092,II3091,WX583);
	nand 	XG13279 	(II3079,II3078,WX582);
	nand 	XG13280 	(II3066,II3065,WX581);
	nand 	XG13281 	(II3053,II3052,WX580);
	nand 	XG13282 	(II3054,II3052,WX485);
	nand 	XG13283 	(II3067,II3065,WX487);
	nand 	XG13284 	(II3080,II3078,WX489);
	nand 	XG13285 	(II3093,II3091,WX491);
	nand 	XG13286 	(II3106,II3104,WX493);
	nand 	XG13287 	(II3119,II3117,WX495);
	nand 	XG13288 	(II3132,II3130,WX497);
	nand 	XG13289 	(II3145,II3143,WX499);
	nand 	XG13290 	(II3158,II3156,WX501);
	nand 	XG13291 	(II3171,II3169,WX503);
	nand 	XG13292 	(II3184,II3182,WX505);
	nand 	XG13293 	(II3197,II3195,WX507);
	nand 	XG13294 	(II3210,II3208,WX509);
	nand 	XG13295 	(II3223,II3221,WX511);
	nand 	XG13296 	(II3236,II3234,WX513);
	nand 	XG13297 	(II3249,II3247,WX515);
	nand 	XG13298 	(II3262,II3260,WX517);
	nand 	XG13299 	(II3275,II3273,WX519);
	nand 	XG13300 	(II3288,II3286,WX521);
	nand 	XG13301 	(II3301,II3299,WX523);
	nand 	XG13302 	(II3314,II3312,WX525);
	nand 	XG13303 	(II3327,II3325,WX527);
	nand 	XG13304 	(II3340,II3338,WX529);
	nand 	XG13305 	(II3353,II3351,WX531);
	nand 	XG13306 	(II3366,II3364,WX533);
	nand 	XG13307 	(II3379,II3377,WX535);
	nand 	XG13308 	(II3392,II3390,WX537);
	nand 	XG13309 	(II3405,II3403,WX539);
	nand 	XG13310 	(II3418,II3416,WX541);
	nand 	XG13311 	(II3431,II3429,WX543);
	nand 	XG13312 	(II3444,II3442,WX545);
	nand 	XG13313 	(II3457,II3455,WX547);
	nand 	XG13314 	(II7059,II7057,WX1778);
	nand 	XG13315 	(II7072,II7070,WX1780);
	nand 	XG13316 	(II7085,II7083,WX1782);
	nand 	XG13317 	(II7098,II7096,WX1784);
	nand 	XG13318 	(II7111,II7109,WX1786);
	nand 	XG13319 	(II7124,II7122,WX1788);
	nand 	XG13320 	(II7137,II7135,WX1790);
	nand 	XG13321 	(II7150,II7148,WX1792);
	nand 	XG13322 	(II7163,II7161,WX1794);
	nand 	XG13323 	(II7176,II7174,WX1796);
	nand 	XG13324 	(II7189,II7187,WX1798);
	nand 	XG13325 	(II7202,II7200,WX1800);
	nand 	XG13326 	(II7215,II7213,WX1802);
	nand 	XG13327 	(II7228,II7226,WX1804);
	nand 	XG13328 	(II7241,II7239,WX1806);
	nand 	XG13329 	(II7254,II7252,WX1808);
	nand 	XG13330 	(II7267,II7265,WX1810);
	nand 	XG13331 	(II7280,II7278,WX1812);
	nand 	XG13332 	(II7293,II7291,WX1814);
	nand 	XG13333 	(II7306,II7304,WX1816);
	nand 	XG13334 	(II7319,II7317,WX1818);
	nand 	XG13335 	(II7332,II7330,WX1820);
	nand 	XG13336 	(II7345,II7343,WX1822);
	nand 	XG13337 	(II7358,II7356,WX1824);
	nand 	XG13338 	(II7371,II7369,WX1826);
	nand 	XG13339 	(II7384,II7382,WX1828);
	nand 	XG13340 	(II7397,II7395,WX1830);
	nand 	XG13341 	(II7410,II7408,WX1832);
	nand 	XG13342 	(II7423,II7421,WX1834);
	nand 	XG13343 	(II7436,II7434,WX1836);
	nand 	XG13344 	(II7449,II7447,WX1838);
	nand 	XG13345 	(II7462,II7460,WX1840);
	nand 	XG13346 	(II11064,II11062,WX3071);
	nand 	XG13347 	(II11077,II11075,WX3073);
	nand 	XG13348 	(II11090,II11088,WX3075);
	nand 	XG13349 	(II11103,II11101,WX3077);
	nand 	XG13350 	(II11116,II11114,WX3079);
	nand 	XG13351 	(II11129,II11127,WX3081);
	nand 	XG13352 	(II11142,II11140,WX3083);
	nand 	XG13353 	(II11155,II11153,WX3085);
	nand 	XG13354 	(II11168,II11166,WX3087);
	nand 	XG13355 	(II11181,II11179,WX3089);
	nand 	XG13356 	(II11194,II11192,WX3091);
	nand 	XG13357 	(II11207,II11205,WX3093);
	nand 	XG13358 	(II11220,II11218,WX3095);
	nand 	XG13359 	(II11233,II11231,WX3097);
	nand 	XG13360 	(II11246,II11244,WX3099);
	nand 	XG13361 	(II11259,II11257,WX3101);
	nand 	XG13362 	(II11272,II11270,WX3103);
	nand 	XG13363 	(II11285,II11283,WX3105);
	nand 	XG13364 	(II11298,II11296,WX3107);
	nand 	XG13365 	(II11311,II11309,WX3109);
	nand 	XG13366 	(II11324,II11322,WX3111);
	nand 	XG13367 	(II11337,II11335,WX3113);
	nand 	XG13368 	(II11350,II11348,WX3115);
	nand 	XG13369 	(II11363,II11361,WX3117);
	nand 	XG13370 	(II11376,II11374,WX3119);
	nand 	XG13371 	(II11389,II11387,WX3121);
	nand 	XG13372 	(II11402,II11400,WX3123);
	nand 	XG13373 	(II11415,II11413,WX3125);
	nand 	XG13374 	(II11428,II11426,WX3127);
	nand 	XG13375 	(II11441,II11439,WX3129);
	nand 	XG13376 	(II11454,II11452,WX3131);
	nand 	XG13377 	(II11467,II11465,WX3133);
	nand 	XG13378 	(II15069,II15067,WX4364);
	nand 	XG13379 	(II15082,II15080,WX4366);
	nand 	XG13380 	(II15095,II15093,WX4368);
	nand 	XG13381 	(II15108,II15106,WX4370);
	nand 	XG13382 	(II15121,II15119,WX4372);
	nand 	XG13383 	(II15134,II15132,WX4374);
	nand 	XG13384 	(II15147,II15145,WX4376);
	nand 	XG13385 	(II15160,II15158,WX4378);
	nand 	XG13386 	(II15173,II15171,WX4380);
	nand 	XG13387 	(II15186,II15184,WX4382);
	nand 	XG13388 	(II15199,II15197,WX4384);
	nand 	XG13389 	(II15212,II15210,WX4386);
	nand 	XG13390 	(II15225,II15223,WX4388);
	nand 	XG13391 	(II15238,II15236,WX4390);
	nand 	XG13392 	(II15251,II15249,WX4392);
	nand 	XG13393 	(II15264,II15262,WX4394);
	nand 	XG13394 	(II15277,II15275,WX4396);
	nand 	XG13395 	(II15290,II15288,WX4398);
	nand 	XG13396 	(II15303,II15301,WX4400);
	nand 	XG13397 	(II15316,II15314,WX4402);
	nand 	XG13398 	(II15329,II15327,WX4404);
	nand 	XG13399 	(II15342,II15340,WX4406);
	nand 	XG13400 	(II15355,II15353,WX4408);
	nand 	XG13401 	(II15368,II15366,WX4410);
	nand 	XG13402 	(II15381,II15379,WX4412);
	nand 	XG13403 	(II15394,II15392,WX4414);
	nand 	XG13404 	(II15407,II15405,WX4416);
	nand 	XG13405 	(II15420,II15418,WX4418);
	nand 	XG13406 	(II15433,II15431,WX4420);
	nand 	XG13407 	(II15446,II15444,WX4422);
	nand 	XG13408 	(II15459,II15457,WX4424);
	nand 	XG13409 	(II15472,II15470,WX4426);
	nand 	XG13410 	(II19074,II19072,WX5657);
	nand 	XG13411 	(II19087,II19085,WX5659);
	nand 	XG13412 	(II19100,II19098,WX5661);
	nand 	XG13413 	(II19113,II19111,WX5663);
	nand 	XG13414 	(II19126,II19124,WX5665);
	nand 	XG13415 	(II19139,II19137,WX5667);
	nand 	XG13416 	(II19152,II19150,WX5669);
	nand 	XG13417 	(II19165,II19163,WX5671);
	nand 	XG13418 	(II19178,II19176,WX5673);
	nand 	XG13419 	(II19191,II19189,WX5675);
	nand 	XG13420 	(II19204,II19202,WX5677);
	nand 	XG13421 	(II19217,II19215,WX5679);
	nand 	XG13422 	(II19230,II19228,WX5681);
	nand 	XG13423 	(II19243,II19241,WX5683);
	nand 	XG13424 	(II19256,II19254,WX5685);
	nand 	XG13425 	(II19269,II19267,WX5687);
	nand 	XG13426 	(II19282,II19280,WX5689);
	nand 	XG13427 	(II19295,II19293,WX5691);
	nand 	XG13428 	(II19308,II19306,WX5693);
	nand 	XG13429 	(II19321,II19319,WX5695);
	nand 	XG13430 	(II19334,II19332,WX5697);
	nand 	XG13431 	(II19347,II19345,WX5699);
	nand 	XG13432 	(II19360,II19358,WX5701);
	nand 	XG13433 	(II19373,II19371,WX5703);
	nand 	XG13434 	(II19386,II19384,WX5705);
	nand 	XG13435 	(II19399,II19397,WX5707);
	nand 	XG13436 	(II19412,II19410,WX5709);
	nand 	XG13437 	(II19425,II19423,WX5711);
	nand 	XG13438 	(II19438,II19436,WX5713);
	nand 	XG13439 	(II19451,II19449,WX5715);
	nand 	XG13440 	(II19464,II19462,WX5717);
	nand 	XG13441 	(II19477,II19475,WX5719);
	nand 	XG13442 	(II23079,II23077,WX6950);
	nand 	XG13443 	(II23092,II23090,WX6952);
	nand 	XG13444 	(II23105,II23103,WX6954);
	nand 	XG13445 	(II23118,II23116,WX6956);
	nand 	XG13446 	(II23131,II23129,WX6958);
	nand 	XG13447 	(II23144,II23142,WX6960);
	nand 	XG13448 	(II23157,II23155,WX6962);
	nand 	XG13449 	(II23170,II23168,WX6964);
	nand 	XG13450 	(II23183,II23181,WX6966);
	nand 	XG13451 	(II23196,II23194,WX6968);
	nand 	XG13452 	(II23209,II23207,WX6970);
	nand 	XG13453 	(II23222,II23220,WX6972);
	nand 	XG13454 	(II23235,II23233,WX6974);
	nand 	XG13455 	(II23248,II23246,WX6976);
	nand 	XG13456 	(II23261,II23259,WX6978);
	nand 	XG13457 	(II23274,II23272,WX6980);
	nand 	XG13458 	(II23287,II23285,WX6982);
	nand 	XG13459 	(II23300,II23298,WX6984);
	nand 	XG13460 	(II23313,II23311,WX6986);
	nand 	XG13461 	(II23326,II23324,WX6988);
	nand 	XG13462 	(II23339,II23337,WX6990);
	nand 	XG13463 	(II23352,II23350,WX6992);
	nand 	XG13464 	(II23365,II23363,WX6994);
	nand 	XG13465 	(II23378,II23376,WX6996);
	nand 	XG13466 	(II23391,II23389,WX6998);
	nand 	XG13467 	(II23404,II23402,WX7000);
	nand 	XG13468 	(II23417,II23415,WX7002);
	nand 	XG13469 	(II23430,II23428,WX7004);
	nand 	XG13470 	(II23443,II23441,WX7006);
	nand 	XG13471 	(II23456,II23454,WX7008);
	nand 	XG13472 	(II23469,II23467,WX7010);
	nand 	XG13473 	(II23482,II23480,WX7012);
	nand 	XG13474 	(II27084,II27082,WX8243);
	nand 	XG13475 	(II27097,II27095,WX8245);
	nand 	XG13476 	(II27110,II27108,WX8247);
	nand 	XG13477 	(II27123,II27121,WX8249);
	nand 	XG13478 	(II27136,II27134,WX8251);
	nand 	XG13479 	(II27149,II27147,WX8253);
	nand 	XG13480 	(II27162,II27160,WX8255);
	nand 	XG13481 	(II27175,II27173,WX8257);
	nand 	XG13482 	(II27188,II27186,WX8259);
	nand 	XG13483 	(II27201,II27199,WX8261);
	nand 	XG13484 	(II27214,II27212,WX8263);
	nand 	XG13485 	(II27227,II27225,WX8265);
	nand 	XG13486 	(II27240,II27238,WX8267);
	nand 	XG13487 	(II27253,II27251,WX8269);
	nand 	XG13488 	(II27266,II27264,WX8271);
	nand 	XG13489 	(II27279,II27277,WX8273);
	nand 	XG13490 	(II27292,II27290,WX8275);
	nand 	XG13491 	(II27305,II27303,WX8277);
	nand 	XG13492 	(II27318,II27316,WX8279);
	nand 	XG13493 	(II27331,II27329,WX8281);
	nand 	XG13494 	(II27344,II27342,WX8283);
	nand 	XG13495 	(II27357,II27355,WX8285);
	nand 	XG13496 	(II27370,II27368,WX8287);
	nand 	XG13497 	(II27383,II27381,WX8289);
	nand 	XG13498 	(II27396,II27394,WX8291);
	nand 	XG13499 	(II27409,II27407,WX8293);
	nand 	XG13500 	(II27422,II27420,WX8295);
	nand 	XG13501 	(II27435,II27433,WX8297);
	nand 	XG13502 	(II27448,II27446,WX8299);
	nand 	XG13503 	(II27461,II27459,WX8301);
	nand 	XG13504 	(II27474,II27472,WX8303);
	nand 	XG13505 	(II27487,II27485,WX8305);
	nand 	XG13506 	(II31089,II31087,WX9536);
	nand 	XG13507 	(II31102,II31100,WX9538);
	nand 	XG13508 	(II31115,II31113,WX9540);
	nand 	XG13509 	(II31128,II31126,WX9542);
	nand 	XG13510 	(II31141,II31139,WX9544);
	nand 	XG13511 	(II31154,II31152,WX9546);
	nand 	XG13512 	(II31167,II31165,WX9548);
	nand 	XG13513 	(II31180,II31178,WX9550);
	nand 	XG13514 	(II31193,II31191,WX9552);
	nand 	XG13515 	(II31206,II31204,WX9554);
	nand 	XG13516 	(II31219,II31217,WX9556);
	nand 	XG13517 	(II31232,II31230,WX9558);
	nand 	XG13518 	(II31245,II31243,WX9560);
	nand 	XG13519 	(II31258,II31256,WX9562);
	nand 	XG13520 	(II31271,II31269,WX9564);
	nand 	XG13521 	(II31284,II31282,WX9566);
	nand 	XG13522 	(II31297,II31295,WX9568);
	nand 	XG13523 	(II31310,II31308,WX9570);
	nand 	XG13524 	(II31323,II31321,WX9572);
	nand 	XG13525 	(II31336,II31334,WX9574);
	nand 	XG13526 	(II31349,II31347,WX9576);
	nand 	XG13527 	(II31362,II31360,WX9578);
	nand 	XG13528 	(II31375,II31373,WX9580);
	nand 	XG13529 	(II31388,II31386,WX9582);
	nand 	XG13530 	(II31401,II31399,WX9584);
	nand 	XG13531 	(II31414,II31412,WX9586);
	nand 	XG13532 	(II31427,II31425,WX9588);
	nand 	XG13533 	(II31440,II31438,WX9590);
	nand 	XG13534 	(II31453,II31451,WX9592);
	nand 	XG13535 	(II31466,II31464,WX9594);
	nand 	XG13536 	(II31479,II31477,WX9596);
	nand 	XG13537 	(II31492,II31490,WX9598);
	nand 	XG13538 	(II35094,II35092,WX10829);
	nand 	XG13539 	(II35107,II35105,WX10831);
	nand 	XG13540 	(II35120,II35118,WX10833);
	nand 	XG13541 	(II35133,II35131,WX10835);
	nand 	XG13542 	(II35146,II35144,WX10837);
	nand 	XG13543 	(II35159,II35157,WX10839);
	nand 	XG13544 	(II35172,II35170,WX10841);
	nand 	XG13545 	(II35185,II35183,WX10843);
	nand 	XG13546 	(II35198,II35196,WX10845);
	nand 	XG13547 	(II35211,II35209,WX10847);
	nand 	XG13548 	(II35224,II35222,WX10849);
	nand 	XG13549 	(II35237,II35235,WX10851);
	nand 	XG13550 	(II35250,II35248,WX10853);
	nand 	XG13551 	(II35263,II35261,WX10855);
	nand 	XG13552 	(II35276,II35274,WX10857);
	nand 	XG13553 	(II35289,II35287,WX10859);
	nand 	XG13554 	(II35302,II35300,WX10861);
	nand 	XG13555 	(II35315,II35313,WX10863);
	nand 	XG13556 	(II35328,II35326,WX10865);
	nand 	XG13557 	(II35341,II35339,WX10867);
	nand 	XG13558 	(II35354,II35352,WX10869);
	nand 	XG13559 	(II35367,II35365,WX10871);
	nand 	XG13560 	(II35380,II35378,WX10873);
	nand 	XG13561 	(II35393,II35391,WX10875);
	nand 	XG13562 	(II35406,II35404,WX10877);
	nand 	XG13563 	(II35419,II35417,WX10879);
	nand 	XG13564 	(II35432,II35430,WX10881);
	nand 	XG13565 	(II35445,II35443,WX10883);
	nand 	XG13566 	(II35458,II35456,WX10885);
	nand 	XG13567 	(II35471,II35469,WX10887);
	nand 	XG13568 	(II35484,II35482,WX10889);
	nand 	XG13569 	(II35497,II35495,WX10891);
	nand 	XG13570 	(WX1006,II3054,II3053);
	nand 	XG13571 	(WX1013,II3067,II3066);
	nand 	XG13572 	(WX1020,II3080,II3079);
	nand 	XG13573 	(WX1027,II3093,II3092);
	nand 	XG13574 	(WX1034,II3106,II3105);
	nand 	XG13575 	(WX1041,II3119,II3118);
	nand 	XG13576 	(WX1048,II3132,II3131);
	nand 	XG13577 	(WX1055,II3145,II3144);
	nand 	XG13578 	(WX1062,II3158,II3157);
	nand 	XG13579 	(WX1069,II3171,II3170);
	nand 	XG13580 	(WX1076,II3184,II3183);
	nand 	XG13581 	(WX1083,II3197,II3196);
	nand 	XG13582 	(WX1090,II3210,II3209);
	nand 	XG13583 	(WX1097,II3223,II3222);
	nand 	XG13584 	(WX1104,II3236,II3235);
	nand 	XG13585 	(WX1111,II3249,II3248);
	nand 	XG13586 	(WX1118,II3262,II3261);
	nand 	XG13587 	(WX1125,II3275,II3274);
	nand 	XG13588 	(WX1132,II3288,II3287);
	nand 	XG13589 	(WX1139,II3301,II3300);
	nand 	XG13590 	(WX1146,II3314,II3313);
	nand 	XG13591 	(WX1153,II3327,II3326);
	nand 	XG13592 	(WX1160,II3340,II3339);
	nand 	XG13593 	(WX1167,II3353,II3352);
	nand 	XG13594 	(WX1174,II3366,II3365);
	nand 	XG13595 	(WX1181,II3379,II3378);
	nand 	XG13596 	(WX1188,II3392,II3391);
	nand 	XG13597 	(WX1195,II3405,II3404);
	nand 	XG13598 	(WX1202,II3418,II3417);
	nand 	XG13599 	(WX1209,II3431,II3430);
	nand 	XG13600 	(WX1216,II3444,II3443);
	nand 	XG13601 	(WX1223,II3457,II3456);
	nand 	XG13602 	(WX2299,II7059,II7058);
	nand 	XG13603 	(WX2306,II7072,II7071);
	nand 	XG13604 	(WX2313,II7085,II7084);
	nand 	XG13605 	(WX2320,II7098,II7097);
	nand 	XG13606 	(WX2327,II7111,II7110);
	nand 	XG13607 	(WX2334,II7124,II7123);
	nand 	XG13608 	(WX2341,II7137,II7136);
	nand 	XG13609 	(WX2348,II7150,II7149);
	nand 	XG13610 	(WX2355,II7163,II7162);
	nand 	XG13611 	(WX2362,II7176,II7175);
	nand 	XG13612 	(WX2369,II7189,II7188);
	nand 	XG13613 	(WX2376,II7202,II7201);
	nand 	XG13614 	(WX2383,II7215,II7214);
	nand 	XG13615 	(WX2390,II7228,II7227);
	nand 	XG13616 	(WX2397,II7241,II7240);
	nand 	XG13617 	(WX2404,II7254,II7253);
	nand 	XG13618 	(WX2411,II7267,II7266);
	nand 	XG13619 	(WX2418,II7280,II7279);
	nand 	XG13620 	(WX2425,II7293,II7292);
	nand 	XG13621 	(WX2432,II7306,II7305);
	nand 	XG13622 	(WX2439,II7319,II7318);
	nand 	XG13623 	(WX2446,II7332,II7331);
	nand 	XG13624 	(WX2453,II7345,II7344);
	nand 	XG13625 	(WX2460,II7358,II7357);
	nand 	XG13626 	(WX2467,II7371,II7370);
	nand 	XG13627 	(WX2474,II7384,II7383);
	nand 	XG13628 	(WX2481,II7397,II7396);
	nand 	XG13629 	(WX2488,II7410,II7409);
	nand 	XG13630 	(WX2495,II7423,II7422);
	nand 	XG13631 	(WX2502,II7436,II7435);
	nand 	XG13632 	(WX2509,II7449,II7448);
	nand 	XG13633 	(WX2516,II7462,II7461);
	nand 	XG13634 	(WX3592,II11064,II11063);
	nand 	XG13635 	(WX3599,II11077,II11076);
	nand 	XG13636 	(WX3606,II11090,II11089);
	nand 	XG13637 	(WX3613,II11103,II11102);
	nand 	XG13638 	(WX3620,II11116,II11115);
	nand 	XG13639 	(WX3627,II11129,II11128);
	nand 	XG13640 	(WX3634,II11142,II11141);
	nand 	XG13641 	(WX3641,II11155,II11154);
	nand 	XG13642 	(WX3648,II11168,II11167);
	nand 	XG13643 	(WX3655,II11181,II11180);
	nand 	XG13644 	(WX3662,II11194,II11193);
	nand 	XG13645 	(WX3669,II11207,II11206);
	nand 	XG13646 	(WX3676,II11220,II11219);
	nand 	XG13647 	(WX3683,II11233,II11232);
	nand 	XG13648 	(WX3690,II11246,II11245);
	nand 	XG13649 	(WX3697,II11259,II11258);
	nand 	XG13650 	(WX3704,II11272,II11271);
	nand 	XG13651 	(WX3711,II11285,II11284);
	nand 	XG13652 	(WX3718,II11298,II11297);
	nand 	XG13653 	(WX3725,II11311,II11310);
	nand 	XG13654 	(WX3732,II11324,II11323);
	nand 	XG13655 	(WX3739,II11337,II11336);
	nand 	XG13656 	(WX3746,II11350,II11349);
	nand 	XG13657 	(WX3753,II11363,II11362);
	nand 	XG13658 	(WX3760,II11376,II11375);
	nand 	XG13659 	(WX3767,II11389,II11388);
	nand 	XG13660 	(WX3774,II11402,II11401);
	nand 	XG13661 	(WX3781,II11415,II11414);
	nand 	XG13662 	(WX3788,II11428,II11427);
	nand 	XG13663 	(WX3795,II11441,II11440);
	nand 	XG13664 	(WX3802,II11454,II11453);
	nand 	XG13665 	(WX3809,II11467,II11466);
	nand 	XG13666 	(WX4885,II15069,II15068);
	nand 	XG13667 	(WX4892,II15082,II15081);
	nand 	XG13668 	(WX4899,II15095,II15094);
	nand 	XG13669 	(WX4906,II15108,II15107);
	nand 	XG13670 	(WX4913,II15121,II15120);
	nand 	XG13671 	(WX4920,II15134,II15133);
	nand 	XG13672 	(WX4927,II15147,II15146);
	nand 	XG13673 	(WX4934,II15160,II15159);
	nand 	XG13674 	(WX4941,II15173,II15172);
	nand 	XG13675 	(WX4948,II15186,II15185);
	nand 	XG13676 	(WX4955,II15199,II15198);
	nand 	XG13677 	(WX4962,II15212,II15211);
	nand 	XG13678 	(WX4969,II15225,II15224);
	nand 	XG13679 	(WX4976,II15238,II15237);
	nand 	XG13680 	(WX4983,II15251,II15250);
	nand 	XG13681 	(WX4990,II15264,II15263);
	nand 	XG13682 	(WX4997,II15277,II15276);
	nand 	XG13683 	(WX5004,II15290,II15289);
	nand 	XG13684 	(WX5011,II15303,II15302);
	nand 	XG13685 	(WX5018,II15316,II15315);
	nand 	XG13686 	(WX5025,II15329,II15328);
	nand 	XG13687 	(WX5032,II15342,II15341);
	nand 	XG13688 	(WX5039,II15355,II15354);
	nand 	XG13689 	(WX5046,II15368,II15367);
	nand 	XG13690 	(WX5053,II15381,II15380);
	nand 	XG13691 	(WX5060,II15394,II15393);
	nand 	XG13692 	(WX5067,II15407,II15406);
	nand 	XG13693 	(WX5074,II15420,II15419);
	nand 	XG13694 	(WX5081,II15433,II15432);
	nand 	XG13695 	(WX5088,II15446,II15445);
	nand 	XG13696 	(WX5095,II15459,II15458);
	nand 	XG13697 	(WX5102,II15472,II15471);
	nand 	XG13698 	(WX6178,II19074,II19073);
	nand 	XG13699 	(WX6185,II19087,II19086);
	nand 	XG13700 	(WX6192,II19100,II19099);
	nand 	XG13701 	(WX6199,II19113,II19112);
	nand 	XG13702 	(WX6206,II19126,II19125);
	nand 	XG13703 	(WX6213,II19139,II19138);
	nand 	XG13704 	(WX6220,II19152,II19151);
	nand 	XG13705 	(WX6227,II19165,II19164);
	nand 	XG13706 	(WX6234,II19178,II19177);
	nand 	XG13707 	(WX6241,II19191,II19190);
	nand 	XG13708 	(WX6248,II19204,II19203);
	nand 	XG13709 	(WX6255,II19217,II19216);
	nand 	XG13710 	(WX6262,II19230,II19229);
	nand 	XG13711 	(WX6269,II19243,II19242);
	nand 	XG13712 	(WX6276,II19256,II19255);
	nand 	XG13713 	(WX6283,II19269,II19268);
	nand 	XG13714 	(WX6290,II19282,II19281);
	nand 	XG13715 	(WX6297,II19295,II19294);
	nand 	XG13716 	(WX6304,II19308,II19307);
	nand 	XG13717 	(WX6311,II19321,II19320);
	nand 	XG13718 	(WX6318,II19334,II19333);
	nand 	XG13719 	(WX6325,II19347,II19346);
	nand 	XG13720 	(WX6332,II19360,II19359);
	nand 	XG13721 	(WX6339,II19373,II19372);
	nand 	XG13722 	(WX6346,II19386,II19385);
	nand 	XG13723 	(WX6353,II19399,II19398);
	nand 	XG13724 	(WX6360,II19412,II19411);
	nand 	XG13725 	(WX6367,II19425,II19424);
	nand 	XG13726 	(WX6374,II19438,II19437);
	nand 	XG13727 	(WX6381,II19451,II19450);
	nand 	XG13728 	(WX6388,II19464,II19463);
	nand 	XG13729 	(WX6395,II19477,II19476);
	nand 	XG13730 	(WX7471,II23079,II23078);
	nand 	XG13731 	(WX7478,II23092,II23091);
	nand 	XG13732 	(WX7485,II23105,II23104);
	nand 	XG13733 	(WX7492,II23118,II23117);
	nand 	XG13734 	(WX7499,II23131,II23130);
	nand 	XG13735 	(WX7506,II23144,II23143);
	nand 	XG13736 	(WX7513,II23157,II23156);
	nand 	XG13737 	(WX7520,II23170,II23169);
	nand 	XG13738 	(WX7527,II23183,II23182);
	nand 	XG13739 	(WX7534,II23196,II23195);
	nand 	XG13740 	(WX7541,II23209,II23208);
	nand 	XG13741 	(WX7548,II23222,II23221);
	nand 	XG13742 	(WX7555,II23235,II23234);
	nand 	XG13743 	(WX7562,II23248,II23247);
	nand 	XG13744 	(WX7569,II23261,II23260);
	nand 	XG13745 	(WX7576,II23274,II23273);
	nand 	XG13746 	(WX7583,II23287,II23286);
	nand 	XG13747 	(WX7590,II23300,II23299);
	nand 	XG13748 	(WX7597,II23313,II23312);
	nand 	XG13749 	(WX7604,II23326,II23325);
	nand 	XG13750 	(WX7611,II23339,II23338);
	nand 	XG13751 	(WX7618,II23352,II23351);
	nand 	XG13752 	(WX7625,II23365,II23364);
	nand 	XG13753 	(WX7632,II23378,II23377);
	nand 	XG13754 	(WX7639,II23391,II23390);
	nand 	XG13755 	(WX7646,II23404,II23403);
	nand 	XG13756 	(WX7653,II23417,II23416);
	nand 	XG13757 	(WX7660,II23430,II23429);
	nand 	XG13758 	(WX7667,II23443,II23442);
	nand 	XG13759 	(WX7674,II23456,II23455);
	nand 	XG13760 	(WX7681,II23469,II23468);
	nand 	XG13761 	(WX7688,II23482,II23481);
	nand 	XG13762 	(WX8764,II27084,II27083);
	nand 	XG13763 	(WX8771,II27097,II27096);
	nand 	XG13764 	(WX8778,II27110,II27109);
	nand 	XG13765 	(WX8785,II27123,II27122);
	nand 	XG13766 	(WX8792,II27136,II27135);
	nand 	XG13767 	(WX8799,II27149,II27148);
	nand 	XG13768 	(WX8806,II27162,II27161);
	nand 	XG13769 	(WX8813,II27175,II27174);
	nand 	XG13770 	(WX8820,II27188,II27187);
	nand 	XG13771 	(WX8827,II27201,II27200);
	nand 	XG13772 	(WX8834,II27214,II27213);
	nand 	XG13773 	(WX8841,II27227,II27226);
	nand 	XG13774 	(WX8848,II27240,II27239);
	nand 	XG13775 	(WX8855,II27253,II27252);
	nand 	XG13776 	(WX8862,II27266,II27265);
	nand 	XG13777 	(WX8869,II27279,II27278);
	nand 	XG13778 	(WX8876,II27292,II27291);
	nand 	XG13779 	(WX8883,II27305,II27304);
	nand 	XG13780 	(WX8890,II27318,II27317);
	nand 	XG13781 	(WX8897,II27331,II27330);
	nand 	XG13782 	(WX8904,II27344,II27343);
	nand 	XG13783 	(WX8911,II27357,II27356);
	nand 	XG13784 	(WX8918,II27370,II27369);
	nand 	XG13785 	(WX8925,II27383,II27382);
	nand 	XG13786 	(WX8932,II27396,II27395);
	nand 	XG13787 	(WX8939,II27409,II27408);
	nand 	XG13788 	(WX8946,II27422,II27421);
	nand 	XG13789 	(WX8953,II27435,II27434);
	nand 	XG13790 	(WX8960,II27448,II27447);
	nand 	XG13791 	(WX8967,II27461,II27460);
	nand 	XG13792 	(WX8974,II27474,II27473);
	nand 	XG13793 	(WX8981,II27487,II27486);
	nand 	XG13794 	(WX10057,II31089,II31088);
	nand 	XG13795 	(WX10064,II31102,II31101);
	nand 	XG13796 	(WX10071,II31115,II31114);
	nand 	XG13797 	(WX10078,II31128,II31127);
	nand 	XG13798 	(WX10085,II31141,II31140);
	nand 	XG13799 	(WX10092,II31154,II31153);
	nand 	XG13800 	(WX10099,II31167,II31166);
	nand 	XG13801 	(WX10106,II31180,II31179);
	nand 	XG13802 	(WX10113,II31193,II31192);
	nand 	XG13803 	(WX10120,II31206,II31205);
	nand 	XG13804 	(WX10127,II31219,II31218);
	nand 	XG13805 	(WX10134,II31232,II31231);
	nand 	XG13806 	(WX10141,II31245,II31244);
	nand 	XG13807 	(WX10148,II31258,II31257);
	nand 	XG13808 	(WX10155,II31271,II31270);
	nand 	XG13809 	(WX10162,II31284,II31283);
	nand 	XG13810 	(WX10169,II31297,II31296);
	nand 	XG13811 	(WX10176,II31310,II31309);
	nand 	XG13812 	(WX10183,II31323,II31322);
	nand 	XG13813 	(WX10190,II31336,II31335);
	nand 	XG13814 	(WX10197,II31349,II31348);
	nand 	XG13815 	(WX10204,II31362,II31361);
	nand 	XG13816 	(WX10211,II31375,II31374);
	nand 	XG13817 	(WX10218,II31388,II31387);
	nand 	XG13818 	(WX10225,II31401,II31400);
	nand 	XG13819 	(WX10232,II31414,II31413);
	nand 	XG13820 	(WX10239,II31427,II31426);
	nand 	XG13821 	(WX10246,II31440,II31439);
	nand 	XG13822 	(WX10253,II31453,II31452);
	nand 	XG13823 	(WX10260,II31466,II31465);
	nand 	XG13824 	(WX10267,II31479,II31478);
	nand 	XG13825 	(WX10274,II31492,II31491);
	nand 	XG13826 	(WX11350,II35094,II35093);
	nand 	XG13827 	(WX11357,II35107,II35106);
	nand 	XG13828 	(WX11364,II35120,II35119);
	nand 	XG13829 	(WX11371,II35133,II35132);
	nand 	XG13830 	(WX11378,II35146,II35145);
	nand 	XG13831 	(WX11385,II35159,II35158);
	nand 	XG13832 	(WX11392,II35172,II35171);
	nand 	XG13833 	(WX11399,II35185,II35184);
	nand 	XG13834 	(WX11406,II35198,II35197);
	nand 	XG13835 	(WX11413,II35211,II35210);
	nand 	XG13836 	(WX11420,II35224,II35223);
	nand 	XG13837 	(WX11427,II35237,II35236);
	nand 	XG13838 	(WX11434,II35250,II35249);
	nand 	XG13839 	(WX11441,II35263,II35262);
	nand 	XG13840 	(WX11448,II35276,II35275);
	nand 	XG13841 	(WX11455,II35289,II35288);
	nand 	XG13842 	(WX11462,II35302,II35301);
	nand 	XG13843 	(WX11469,II35315,II35314);
	nand 	XG13844 	(WX11476,II35328,II35327);
	nand 	XG13845 	(WX11483,II35341,II35340);
	nand 	XG13846 	(WX11490,II35354,II35353);
	nand 	XG13847 	(WX11497,II35367,II35366);
	nand 	XG13848 	(WX11504,II35380,II35379);
	nand 	XG13849 	(WX11511,II35393,II35392);
	nand 	XG13850 	(WX11518,II35406,II35405);
	nand 	XG13851 	(WX11525,II35419,II35418);
	nand 	XG13852 	(WX11532,II35432,II35431);
	nand 	XG13853 	(WX11539,II35445,II35444);
	nand 	XG13854 	(WX11546,II35458,II35457);
	nand 	XG13855 	(WX11553,II35471,II35470);
	nand 	XG13856 	(WX11560,II35484,II35483);
	nand 	XG13857 	(WX11567,II35497,II35496);
	and 	XG13858 	(WX11568,WX11349,WX11567);
	and 	XG13859 	(WX11561,WX11349,WX11560);
	and 	XG13860 	(WX11554,WX11349,WX11553);
	and 	XG13861 	(WX11547,WX11349,WX11546);
	and 	XG13862 	(WX11540,WX11349,WX11539);
	and 	XG13863 	(WX11533,WX11349,WX11532);
	and 	XG13864 	(WX11526,WX11349,WX11525);
	and 	XG13865 	(WX11519,WX11349,WX11518);
	and 	XG13866 	(WX11512,WX11349,WX11511);
	and 	XG13867 	(WX11505,WX11349,WX11504);
	and 	XG13868 	(WX11498,WX11349,WX11497);
	and 	XG13869 	(WX11491,WX11349,WX11490);
	and 	XG13870 	(WX11484,WX11349,WX11483);
	and 	XG13871 	(WX11477,WX11349,WX11476);
	and 	XG13872 	(WX11470,WX11349,WX11469);
	and 	XG13873 	(WX11463,WX11349,WX11462);
	and 	XG13874 	(WX11456,WX11349,WX11455);
	and 	XG13875 	(WX11449,WX11349,WX11448);
	and 	XG13876 	(WX11442,WX11349,WX11441);
	and 	XG13877 	(WX11435,WX11349,WX11434);
	and 	XG13878 	(WX11428,WX11349,WX11427);
	and 	XG13879 	(WX11421,WX11349,WX11420);
	and 	XG13880 	(WX11414,WX11349,WX11413);
	and 	XG13881 	(WX11407,WX11349,WX11406);
	and 	XG13882 	(WX11400,WX11349,WX11399);
	and 	XG13883 	(WX11393,WX11349,WX11392);
	and 	XG13884 	(WX11386,WX11349,WX11385);
	and 	XG13885 	(WX11379,WX11349,WX11378);
	and 	XG13886 	(WX11372,WX11349,WX11371);
	and 	XG13887 	(WX11365,WX11349,WX11364);
	and 	XG13888 	(WX11358,WX11349,WX11357);
	and 	XG13889 	(WX11351,WX11349,WX11350);
	and 	XG13890 	(WX10275,WX10056,WX10274);
	and 	XG13891 	(WX10268,WX10056,WX10267);
	and 	XG13892 	(WX10261,WX10056,WX10260);
	and 	XG13893 	(WX10254,WX10056,WX10253);
	and 	XG13894 	(WX10247,WX10056,WX10246);
	and 	XG13895 	(WX10240,WX10056,WX10239);
	and 	XG13896 	(WX10233,WX10056,WX10232);
	and 	XG13897 	(WX10226,WX10056,WX10225);
	and 	XG13898 	(WX10219,WX10056,WX10218);
	and 	XG13899 	(WX10212,WX10056,WX10211);
	and 	XG13900 	(WX10205,WX10056,WX10204);
	and 	XG13901 	(WX10198,WX10056,WX10197);
	and 	XG13902 	(WX10191,WX10056,WX10190);
	and 	XG13903 	(WX10184,WX10056,WX10183);
	and 	XG13904 	(WX10177,WX10056,WX10176);
	and 	XG13905 	(WX10170,WX10056,WX10169);
	and 	XG13906 	(WX10163,WX10056,WX10162);
	and 	XG13907 	(WX10156,WX10056,WX10155);
	and 	XG13908 	(WX10149,WX10056,WX10148);
	and 	XG13909 	(WX10142,WX10056,WX10141);
	and 	XG13910 	(WX10135,WX10056,WX10134);
	and 	XG13911 	(WX10128,WX10056,WX10127);
	and 	XG13912 	(WX10121,WX10056,WX10120);
	and 	XG13913 	(WX10114,WX10056,WX10113);
	and 	XG13914 	(WX10107,WX10056,WX10106);
	and 	XG13915 	(WX10100,WX10056,WX10099);
	and 	XG13916 	(WX10093,WX10056,WX10092);
	and 	XG13917 	(WX10086,WX10056,WX10085);
	and 	XG13918 	(WX10079,WX10056,WX10078);
	and 	XG13919 	(WX10072,WX10056,WX10071);
	and 	XG13920 	(WX10065,WX10056,WX10064);
	and 	XG13921 	(WX10058,WX10056,WX10057);
	and 	XG13922 	(WX8982,WX8763,WX8981);
	and 	XG13923 	(WX8975,WX8763,WX8974);
	and 	XG13924 	(WX8968,WX8763,WX8967);
	and 	XG13925 	(WX8961,WX8763,WX8960);
	and 	XG13926 	(WX8954,WX8763,WX8953);
	and 	XG13927 	(WX8947,WX8763,WX8946);
	and 	XG13928 	(WX8940,WX8763,WX8939);
	and 	XG13929 	(WX8933,WX8763,WX8932);
	and 	XG13930 	(WX8926,WX8763,WX8925);
	and 	XG13931 	(WX8919,WX8763,WX8918);
	and 	XG13932 	(WX8912,WX8763,WX8911);
	and 	XG13933 	(WX8905,WX8763,WX8904);
	and 	XG13934 	(WX8898,WX8763,WX8897);
	and 	XG13935 	(WX8891,WX8763,WX8890);
	and 	XG13936 	(WX8884,WX8763,WX8883);
	and 	XG13937 	(WX8877,WX8763,WX8876);
	and 	XG13938 	(WX8870,WX8763,WX8869);
	and 	XG13939 	(WX8863,WX8763,WX8862);
	and 	XG13940 	(WX8856,WX8763,WX8855);
	and 	XG13941 	(WX8849,WX8763,WX8848);
	and 	XG13942 	(WX8842,WX8763,WX8841);
	and 	XG13943 	(WX8835,WX8763,WX8834);
	and 	XG13944 	(WX8828,WX8763,WX8827);
	and 	XG13945 	(WX8821,WX8763,WX8820);
	and 	XG13946 	(WX8814,WX8763,WX8813);
	and 	XG13947 	(WX8807,WX8763,WX8806);
	and 	XG13948 	(WX8800,WX8763,WX8799);
	and 	XG13949 	(WX8793,WX8763,WX8792);
	and 	XG13950 	(WX8786,WX8763,WX8785);
	and 	XG13951 	(WX8779,WX8763,WX8778);
	and 	XG13952 	(WX8772,WX8763,WX8771);
	and 	XG13953 	(WX8765,WX8763,WX8764);
	and 	XG13954 	(WX7689,WX7470,WX7688);
	and 	XG13955 	(WX7682,WX7470,WX7681);
	and 	XG13956 	(WX7675,WX7470,WX7674);
	and 	XG13957 	(WX7668,WX7470,WX7667);
	and 	XG13958 	(WX7661,WX7470,WX7660);
	and 	XG13959 	(WX7654,WX7470,WX7653);
	and 	XG13960 	(WX7647,WX7470,WX7646);
	and 	XG13961 	(WX7640,WX7470,WX7639);
	and 	XG13962 	(WX7633,WX7470,WX7632);
	and 	XG13963 	(WX7626,WX7470,WX7625);
	and 	XG13964 	(WX7619,WX7470,WX7618);
	and 	XG13965 	(WX7612,WX7470,WX7611);
	and 	XG13966 	(WX7605,WX7470,WX7604);
	and 	XG13967 	(WX7598,WX7470,WX7597);
	and 	XG13968 	(WX7591,WX7470,WX7590);
	and 	XG13969 	(WX7584,WX7470,WX7583);
	and 	XG13970 	(WX7577,WX7470,WX7576);
	and 	XG13971 	(WX7570,WX7470,WX7569);
	and 	XG13972 	(WX7563,WX7470,WX7562);
	and 	XG13973 	(WX7556,WX7470,WX7555);
	and 	XG13974 	(WX7549,WX7470,WX7548);
	and 	XG13975 	(WX7542,WX7470,WX7541);
	and 	XG13976 	(WX7535,WX7470,WX7534);
	and 	XG13977 	(WX7528,WX7470,WX7527);
	and 	XG13978 	(WX7521,WX7470,WX7520);
	and 	XG13979 	(WX7514,WX7470,WX7513);
	and 	XG13980 	(WX7507,WX7470,WX7506);
	and 	XG13981 	(WX7500,WX7470,WX7499);
	and 	XG13982 	(WX7493,WX7470,WX7492);
	and 	XG13983 	(WX7486,WX7470,WX7485);
	and 	XG13984 	(WX7479,WX7470,WX7478);
	and 	XG13985 	(WX7472,WX7470,WX7471);
	and 	XG13986 	(WX6396,WX6177,WX6395);
	and 	XG13987 	(WX6389,WX6177,WX6388);
	and 	XG13988 	(WX6382,WX6177,WX6381);
	and 	XG13989 	(WX6375,WX6177,WX6374);
	and 	XG13990 	(WX6368,WX6177,WX6367);
	and 	XG13991 	(WX6361,WX6177,WX6360);
	and 	XG13992 	(WX6354,WX6177,WX6353);
	and 	XG13993 	(WX6347,WX6177,WX6346);
	and 	XG13994 	(WX6340,WX6177,WX6339);
	and 	XG13995 	(WX6333,WX6177,WX6332);
	and 	XG13996 	(WX6326,WX6177,WX6325);
	and 	XG13997 	(WX6319,WX6177,WX6318);
	and 	XG13998 	(WX6312,WX6177,WX6311);
	and 	XG13999 	(WX6305,WX6177,WX6304);
	and 	XG14000 	(WX6298,WX6177,WX6297);
	and 	XG14001 	(WX6291,WX6177,WX6290);
	and 	XG14002 	(WX6284,WX6177,WX6283);
	and 	XG14003 	(WX6277,WX6177,WX6276);
	and 	XG14004 	(WX6270,WX6177,WX6269);
	and 	XG14005 	(WX6263,WX6177,WX6262);
	and 	XG14006 	(WX6256,WX6177,WX6255);
	and 	XG14007 	(WX6249,WX6177,WX6248);
	and 	XG14008 	(WX6242,WX6177,WX6241);
	and 	XG14009 	(WX6235,WX6177,WX6234);
	and 	XG14010 	(WX6228,WX6177,WX6227);
	and 	XG14011 	(WX6221,WX6177,WX6220);
	and 	XG14012 	(WX6214,WX6177,WX6213);
	and 	XG14013 	(WX6207,WX6177,WX6206);
	and 	XG14014 	(WX6200,WX6177,WX6199);
	and 	XG14015 	(WX6193,WX6177,WX6192);
	and 	XG14016 	(WX6186,WX6177,WX6185);
	and 	XG14017 	(WX6179,WX6177,WX6178);
	and 	XG14018 	(WX5103,WX4884,WX5102);
	and 	XG14019 	(WX5096,WX4884,WX5095);
	and 	XG14020 	(WX5089,WX4884,WX5088);
	and 	XG14021 	(WX5082,WX4884,WX5081);
	and 	XG14022 	(WX5075,WX4884,WX5074);
	and 	XG14023 	(WX5068,WX4884,WX5067);
	and 	XG14024 	(WX5061,WX4884,WX5060);
	and 	XG14025 	(WX5054,WX4884,WX5053);
	and 	XG14026 	(WX5047,WX4884,WX5046);
	and 	XG14027 	(WX5040,WX4884,WX5039);
	and 	XG14028 	(WX5033,WX4884,WX5032);
	and 	XG14029 	(WX5026,WX4884,WX5025);
	and 	XG14030 	(WX5019,WX4884,WX5018);
	and 	XG14031 	(WX5012,WX4884,WX5011);
	and 	XG14032 	(WX5005,WX4884,WX5004);
	and 	XG14033 	(WX4998,WX4884,WX4997);
	and 	XG14034 	(WX4991,WX4884,WX4990);
	and 	XG14035 	(WX4984,WX4884,WX4983);
	and 	XG14036 	(WX4977,WX4884,WX4976);
	and 	XG14037 	(WX4970,WX4884,WX4969);
	and 	XG14038 	(WX4963,WX4884,WX4962);
	and 	XG14039 	(WX4956,WX4884,WX4955);
	and 	XG14040 	(WX4949,WX4884,WX4948);
	and 	XG14041 	(WX4942,WX4884,WX4941);
	and 	XG14042 	(WX4935,WX4884,WX4934);
	and 	XG14043 	(WX4928,WX4884,WX4927);
	and 	XG14044 	(WX4921,WX4884,WX4920);
	and 	XG14045 	(WX4914,WX4884,WX4913);
	and 	XG14046 	(WX4907,WX4884,WX4906);
	and 	XG14047 	(WX4900,WX4884,WX4899);
	and 	XG14048 	(WX4893,WX4884,WX4892);
	and 	XG14049 	(WX4886,WX4884,WX4885);
	and 	XG14050 	(WX3810,WX3591,WX3809);
	and 	XG14051 	(WX3803,WX3591,WX3802);
	and 	XG14052 	(WX3796,WX3591,WX3795);
	and 	XG14053 	(WX3789,WX3591,WX3788);
	and 	XG14054 	(WX3782,WX3591,WX3781);
	and 	XG14055 	(WX3775,WX3591,WX3774);
	and 	XG14056 	(WX3768,WX3591,WX3767);
	and 	XG14057 	(WX3761,WX3591,WX3760);
	and 	XG14058 	(WX3754,WX3591,WX3753);
	and 	XG14059 	(WX3747,WX3591,WX3746);
	and 	XG14060 	(WX3740,WX3591,WX3739);
	and 	XG14061 	(WX3733,WX3591,WX3732);
	and 	XG14062 	(WX3726,WX3591,WX3725);
	and 	XG14063 	(WX3719,WX3591,WX3718);
	and 	XG14064 	(WX3712,WX3591,WX3711);
	and 	XG14065 	(WX3705,WX3591,WX3704);
	and 	XG14066 	(WX3698,WX3591,WX3697);
	and 	XG14067 	(WX3691,WX3591,WX3690);
	and 	XG14068 	(WX3684,WX3591,WX3683);
	and 	XG14069 	(WX3677,WX3591,WX3676);
	and 	XG14070 	(WX3670,WX3591,WX3669);
	and 	XG14071 	(WX3663,WX3591,WX3662);
	and 	XG14072 	(WX3656,WX3591,WX3655);
	and 	XG14073 	(WX3649,WX3591,WX3648);
	and 	XG14074 	(WX3642,WX3591,WX3641);
	and 	XG14075 	(WX3635,WX3591,WX3634);
	and 	XG14076 	(WX3628,WX3591,WX3627);
	and 	XG14077 	(WX3621,WX3591,WX3620);
	and 	XG14078 	(WX3614,WX3591,WX3613);
	and 	XG14079 	(WX3607,WX3591,WX3606);
	and 	XG14080 	(WX3600,WX3591,WX3599);
	and 	XG14081 	(WX3593,WX3591,WX3592);
	and 	XG14082 	(WX2517,WX2298,WX2516);
	and 	XG14083 	(WX2510,WX2298,WX2509);
	and 	XG14084 	(WX2503,WX2298,WX2502);
	and 	XG14085 	(WX2496,WX2298,WX2495);
	and 	XG14086 	(WX2489,WX2298,WX2488);
	and 	XG14087 	(WX2482,WX2298,WX2481);
	and 	XG14088 	(WX2475,WX2298,WX2474);
	and 	XG14089 	(WX2468,WX2298,WX2467);
	and 	XG14090 	(WX2461,WX2298,WX2460);
	and 	XG14091 	(WX2454,WX2298,WX2453);
	and 	XG14092 	(WX2447,WX2298,WX2446);
	and 	XG14093 	(WX2440,WX2298,WX2439);
	and 	XG14094 	(WX2433,WX2298,WX2432);
	and 	XG14095 	(WX2426,WX2298,WX2425);
	and 	XG14096 	(WX2419,WX2298,WX2418);
	and 	XG14097 	(WX2412,WX2298,WX2411);
	and 	XG14098 	(WX2405,WX2298,WX2404);
	and 	XG14099 	(WX2398,WX2298,WX2397);
	and 	XG14100 	(WX2391,WX2298,WX2390);
	and 	XG14101 	(WX2384,WX2298,WX2383);
	and 	XG14102 	(WX2377,WX2298,WX2376);
	and 	XG14103 	(WX2370,WX2298,WX2369);
	and 	XG14104 	(WX2363,WX2298,WX2362);
	and 	XG14105 	(WX2356,WX2298,WX2355);
	and 	XG14106 	(WX2349,WX2298,WX2348);
	and 	XG14107 	(WX2342,WX2298,WX2341);
	and 	XG14108 	(WX2335,WX2298,WX2334);
	and 	XG14109 	(WX2328,WX2298,WX2327);
	and 	XG14110 	(WX2321,WX2298,WX2320);
	and 	XG14111 	(WX2314,WX2298,WX2313);
	and 	XG14112 	(WX2307,WX2298,WX2306);
	and 	XG14113 	(WX2300,WX2298,WX2299);
	and 	XG14114 	(WX1224,WX1005,WX1223);
	and 	XG14115 	(WX1217,WX1005,WX1216);
	and 	XG14116 	(WX1210,WX1005,WX1209);
	and 	XG14117 	(WX1203,WX1005,WX1202);
	and 	XG14118 	(WX1196,WX1005,WX1195);
	and 	XG14119 	(WX1189,WX1005,WX1188);
	and 	XG14120 	(WX1182,WX1005,WX1181);
	and 	XG14121 	(WX1175,WX1005,WX1174);
	and 	XG14122 	(WX1168,WX1005,WX1167);
	and 	XG14123 	(WX1161,WX1005,WX1160);
	and 	XG14124 	(WX1154,WX1005,WX1153);
	and 	XG14125 	(WX1147,WX1005,WX1146);
	and 	XG14126 	(WX1140,WX1005,WX1139);
	and 	XG14127 	(WX1133,WX1005,WX1132);
	and 	XG14128 	(WX1126,WX1005,WX1125);
	and 	XG14129 	(WX1119,WX1005,WX1118);
	and 	XG14130 	(WX1112,WX1005,WX1111);
	and 	XG14131 	(WX1105,WX1005,WX1104);
	and 	XG14132 	(WX1098,WX1005,WX1097);
	and 	XG14133 	(WX1091,WX1005,WX1090);
	and 	XG14134 	(WX1084,WX1005,WX1083);
	and 	XG14135 	(WX1077,WX1005,WX1076);
	and 	XG14136 	(WX1070,WX1005,WX1069);
	and 	XG14137 	(WX1063,WX1005,WX1062);
	and 	XG14138 	(WX1056,WX1005,WX1055);
	and 	XG14139 	(WX1049,WX1005,WX1048);
	and 	XG14140 	(WX1042,WX1005,WX1041);
	and 	XG14141 	(WX1035,WX1005,WX1034);
	and 	XG14142 	(WX1028,WX1005,WX1027);
	and 	XG14143 	(WX1021,WX1005,WX1020);
	and 	XG14144 	(WX1014,WX1005,WX1013);
	and 	XG14145 	(WX1007,WX1005,WX1006);
	or 	XG14146 	(WX1010,WX1007,WX1008);
	or 	XG14147 	(WX1017,WX1014,WX1015);
	or 	XG14148 	(WX1024,WX1021,WX1022);
	or 	XG14149 	(WX1031,WX1028,WX1029);
	or 	XG14150 	(WX1038,WX1035,WX1036);
	or 	XG14151 	(WX1045,WX1042,WX1043);
	or 	XG14152 	(WX1052,WX1049,WX1050);
	or 	XG14153 	(WX1059,WX1056,WX1057);
	or 	XG14154 	(WX1066,WX1063,WX1064);
	or 	XG14155 	(WX1073,WX1070,WX1071);
	or 	XG14156 	(WX1080,WX1077,WX1078);
	or 	XG14157 	(WX1087,WX1084,WX1085);
	or 	XG14158 	(WX1094,WX1091,WX1092);
	or 	XG14159 	(WX1101,WX1098,WX1099);
	or 	XG14160 	(WX1108,WX1105,WX1106);
	or 	XG14161 	(WX1115,WX1112,WX1113);
	or 	XG14162 	(WX1122,WX1119,WX1120);
	or 	XG14163 	(WX1129,WX1126,WX1127);
	or 	XG14164 	(WX1136,WX1133,WX1134);
	or 	XG14165 	(WX1143,WX1140,WX1141);
	or 	XG14166 	(WX1150,WX1147,WX1148);
	or 	XG14167 	(WX1157,WX1154,WX1155);
	or 	XG14168 	(WX1164,WX1161,WX1162);
	or 	XG14169 	(WX1171,WX1168,WX1169);
	or 	XG14170 	(WX1178,WX1175,WX1176);
	or 	XG14171 	(WX1185,WX1182,WX1183);
	or 	XG14172 	(WX1192,WX1189,WX1190);
	or 	XG14173 	(WX1199,WX1196,WX1197);
	or 	XG14174 	(WX1206,WX1203,WX1204);
	or 	XG14175 	(WX1213,WX1210,WX1211);
	or 	XG14176 	(WX1220,WX1217,WX1218);
	or 	XG14177 	(WX1227,WX1224,WX1225);
	or 	XG14178 	(WX2303,WX2300,WX2301);
	or 	XG14179 	(WX2310,WX2307,WX2308);
	or 	XG14180 	(WX2317,WX2314,WX2315);
	or 	XG14181 	(WX2324,WX2321,WX2322);
	or 	XG14182 	(WX2331,WX2328,WX2329);
	or 	XG14183 	(WX2338,WX2335,WX2336);
	or 	XG14184 	(WX2345,WX2342,WX2343);
	or 	XG14185 	(WX2352,WX2349,WX2350);
	or 	XG14186 	(WX2359,WX2356,WX2357);
	or 	XG14187 	(WX2366,WX2363,WX2364);
	or 	XG14188 	(WX2373,WX2370,WX2371);
	or 	XG14189 	(WX2380,WX2377,WX2378);
	or 	XG14190 	(WX2387,WX2384,WX2385);
	or 	XG14191 	(WX2394,WX2391,WX2392);
	or 	XG14192 	(WX2401,WX2398,WX2399);
	or 	XG14193 	(WX2408,WX2405,WX2406);
	or 	XG14194 	(WX2415,WX2412,WX2413);
	or 	XG14195 	(WX2422,WX2419,WX2420);
	or 	XG14196 	(WX2429,WX2426,WX2427);
	or 	XG14197 	(WX2436,WX2433,WX2434);
	or 	XG14198 	(WX2443,WX2440,WX2441);
	or 	XG14199 	(WX2450,WX2447,WX2448);
	or 	XG14200 	(WX2457,WX2454,WX2455);
	or 	XG14201 	(WX2464,WX2461,WX2462);
	or 	XG14202 	(WX2471,WX2468,WX2469);
	or 	XG14203 	(WX2478,WX2475,WX2476);
	or 	XG14204 	(WX2485,WX2482,WX2483);
	or 	XG14205 	(WX2492,WX2489,WX2490);
	or 	XG14206 	(WX2499,WX2496,WX2497);
	or 	XG14207 	(WX2506,WX2503,WX2504);
	or 	XG14208 	(WX2513,WX2510,WX2511);
	or 	XG14209 	(WX2520,WX2517,WX2518);
	or 	XG14210 	(WX3596,WX3593,WX3594);
	or 	XG14211 	(WX3603,WX3600,WX3601);
	or 	XG14212 	(WX3610,WX3607,WX3608);
	or 	XG14213 	(WX3617,WX3614,WX3615);
	or 	XG14214 	(WX3624,WX3621,WX3622);
	or 	XG14215 	(WX3631,WX3628,WX3629);
	or 	XG14216 	(WX3638,WX3635,WX3636);
	or 	XG14217 	(WX3645,WX3642,WX3643);
	or 	XG14218 	(WX3652,WX3649,WX3650);
	or 	XG14219 	(WX3659,WX3656,WX3657);
	or 	XG14220 	(WX3666,WX3663,WX3664);
	or 	XG14221 	(WX3673,WX3670,WX3671);
	or 	XG14222 	(WX3680,WX3677,WX3678);
	or 	XG14223 	(WX3687,WX3684,WX3685);
	or 	XG14224 	(WX3694,WX3691,WX3692);
	or 	XG14225 	(WX3701,WX3698,WX3699);
	or 	XG14226 	(WX3708,WX3705,WX3706);
	or 	XG14227 	(WX3715,WX3712,WX3713);
	or 	XG14228 	(WX3722,WX3719,WX3720);
	or 	XG14229 	(WX3729,WX3726,WX3727);
	or 	XG14230 	(WX3736,WX3733,WX3734);
	or 	XG14231 	(WX3743,WX3740,WX3741);
	or 	XG14232 	(WX3750,WX3747,WX3748);
	or 	XG14233 	(WX3757,WX3754,WX3755);
	or 	XG14234 	(WX3764,WX3761,WX3762);
	or 	XG14235 	(WX3771,WX3768,WX3769);
	or 	XG14236 	(WX3778,WX3775,WX3776);
	or 	XG14237 	(WX3785,WX3782,WX3783);
	or 	XG14238 	(WX3792,WX3789,WX3790);
	or 	XG14239 	(WX3799,WX3796,WX3797);
	or 	XG14240 	(WX3806,WX3803,WX3804);
	or 	XG14241 	(WX3813,WX3810,WX3811);
	or 	XG14242 	(WX4889,WX4886,WX4887);
	or 	XG14243 	(WX4896,WX4893,WX4894);
	or 	XG14244 	(WX4903,WX4900,WX4901);
	or 	XG14245 	(WX4910,WX4907,WX4908);
	or 	XG14246 	(WX4917,WX4914,WX4915);
	or 	XG14247 	(WX4924,WX4921,WX4922);
	or 	XG14248 	(WX4931,WX4928,WX4929);
	or 	XG14249 	(WX4938,WX4935,WX4936);
	or 	XG14250 	(WX4945,WX4942,WX4943);
	or 	XG14251 	(WX4952,WX4949,WX4950);
	or 	XG14252 	(WX4959,WX4956,WX4957);
	or 	XG14253 	(WX4966,WX4963,WX4964);
	or 	XG14254 	(WX4973,WX4970,WX4971);
	or 	XG14255 	(WX4980,WX4977,WX4978);
	or 	XG14256 	(WX4987,WX4984,WX4985);
	or 	XG14257 	(WX4994,WX4991,WX4992);
	or 	XG14258 	(WX5001,WX4998,WX4999);
	or 	XG14259 	(WX5008,WX5005,WX5006);
	or 	XG14260 	(WX5015,WX5012,WX5013);
	or 	XG14261 	(WX5022,WX5019,WX5020);
	or 	XG14262 	(WX5029,WX5026,WX5027);
	or 	XG14263 	(WX5036,WX5033,WX5034);
	or 	XG14264 	(WX5043,WX5040,WX5041);
	or 	XG14265 	(WX5050,WX5047,WX5048);
	or 	XG14266 	(WX5057,WX5054,WX5055);
	or 	XG14267 	(WX5064,WX5061,WX5062);
	or 	XG14268 	(WX5071,WX5068,WX5069);
	or 	XG14269 	(WX5078,WX5075,WX5076);
	or 	XG14270 	(WX5085,WX5082,WX5083);
	or 	XG14271 	(WX5092,WX5089,WX5090);
	or 	XG14272 	(WX5099,WX5096,WX5097);
	or 	XG14273 	(WX5106,WX5103,WX5104);
	or 	XG14274 	(WX6182,WX6179,WX6180);
	or 	XG14275 	(WX6189,WX6186,WX6187);
	or 	XG14276 	(WX6196,WX6193,WX6194);
	or 	XG14277 	(WX6203,WX6200,WX6201);
	or 	XG14278 	(WX6210,WX6207,WX6208);
	or 	XG14279 	(WX6217,WX6214,WX6215);
	or 	XG14280 	(WX6224,WX6221,WX6222);
	or 	XG14281 	(WX6231,WX6228,WX6229);
	or 	XG14282 	(WX6238,WX6235,WX6236);
	or 	XG14283 	(WX6245,WX6242,WX6243);
	or 	XG14284 	(WX6252,WX6249,WX6250);
	or 	XG14285 	(WX6259,WX6256,WX6257);
	or 	XG14286 	(WX6266,WX6263,WX6264);
	or 	XG14287 	(WX6273,WX6270,WX6271);
	or 	XG14288 	(WX6280,WX6277,WX6278);
	or 	XG14289 	(WX6287,WX6284,WX6285);
	or 	XG14290 	(WX6294,WX6291,WX6292);
	or 	XG14291 	(WX6301,WX6298,WX6299);
	or 	XG14292 	(WX6308,WX6305,WX6306);
	or 	XG14293 	(WX6315,WX6312,WX6313);
	or 	XG14294 	(WX6322,WX6319,WX6320);
	or 	XG14295 	(WX6329,WX6326,WX6327);
	or 	XG14296 	(WX6336,WX6333,WX6334);
	or 	XG14297 	(WX6343,WX6340,WX6341);
	or 	XG14298 	(WX6350,WX6347,WX6348);
	or 	XG14299 	(WX6357,WX6354,WX6355);
	or 	XG14300 	(WX6364,WX6361,WX6362);
	or 	XG14301 	(WX6371,WX6368,WX6369);
	or 	XG14302 	(WX6378,WX6375,WX6376);
	or 	XG14303 	(WX6385,WX6382,WX6383);
	or 	XG14304 	(WX6392,WX6389,WX6390);
	or 	XG14305 	(WX6399,WX6396,WX6397);
	or 	XG14306 	(WX7475,WX7472,WX7473);
	or 	XG14307 	(WX7482,WX7479,WX7480);
	or 	XG14308 	(WX7489,WX7486,WX7487);
	or 	XG14309 	(WX7496,WX7493,WX7494);
	or 	XG14310 	(WX7503,WX7500,WX7501);
	or 	XG14311 	(WX7510,WX7507,WX7508);
	or 	XG14312 	(WX7517,WX7514,WX7515);
	or 	XG14313 	(WX7524,WX7521,WX7522);
	or 	XG14314 	(WX7531,WX7528,WX7529);
	or 	XG14315 	(WX7538,WX7535,WX7536);
	or 	XG14316 	(WX7545,WX7542,WX7543);
	or 	XG14317 	(WX7552,WX7549,WX7550);
	or 	XG14318 	(WX7559,WX7556,WX7557);
	or 	XG14319 	(WX7566,WX7563,WX7564);
	or 	XG14320 	(WX7573,WX7570,WX7571);
	or 	XG14321 	(WX7580,WX7577,WX7578);
	or 	XG14322 	(WX7587,WX7584,WX7585);
	or 	XG14323 	(WX7594,WX7591,WX7592);
	or 	XG14324 	(WX7601,WX7598,WX7599);
	or 	XG14325 	(WX7608,WX7605,WX7606);
	or 	XG14326 	(WX7615,WX7612,WX7613);
	or 	XG14327 	(WX7622,WX7619,WX7620);
	or 	XG14328 	(WX7629,WX7626,WX7627);
	or 	XG14329 	(WX7636,WX7633,WX7634);
	or 	XG14330 	(WX7643,WX7640,WX7641);
	or 	XG14331 	(WX7650,WX7647,WX7648);
	or 	XG14332 	(WX7657,WX7654,WX7655);
	or 	XG14333 	(WX7664,WX7661,WX7662);
	or 	XG14334 	(WX7671,WX7668,WX7669);
	or 	XG14335 	(WX7678,WX7675,WX7676);
	or 	XG14336 	(WX7685,WX7682,WX7683);
	or 	XG14337 	(WX7692,WX7689,WX7690);
	or 	XG14338 	(WX8768,WX8765,WX8766);
	or 	XG14339 	(WX8775,WX8772,WX8773);
	or 	XG14340 	(WX8782,WX8779,WX8780);
	or 	XG14341 	(WX8789,WX8786,WX8787);
	or 	XG14342 	(WX8796,WX8793,WX8794);
	or 	XG14343 	(WX8803,WX8800,WX8801);
	or 	XG14344 	(WX8810,WX8807,WX8808);
	or 	XG14345 	(WX8817,WX8814,WX8815);
	or 	XG14346 	(WX8824,WX8821,WX8822);
	or 	XG14347 	(WX8831,WX8828,WX8829);
	or 	XG14348 	(WX8838,WX8835,WX8836);
	or 	XG14349 	(WX8845,WX8842,WX8843);
	or 	XG14350 	(WX8852,WX8849,WX8850);
	or 	XG14351 	(WX8859,WX8856,WX8857);
	or 	XG14352 	(WX8866,WX8863,WX8864);
	or 	XG14353 	(WX8873,WX8870,WX8871);
	or 	XG14354 	(WX8880,WX8877,WX8878);
	or 	XG14355 	(WX8887,WX8884,WX8885);
	or 	XG14356 	(WX8894,WX8891,WX8892);
	or 	XG14357 	(WX8901,WX8898,WX8899);
	or 	XG14358 	(WX8908,WX8905,WX8906);
	or 	XG14359 	(WX8915,WX8912,WX8913);
	or 	XG14360 	(WX8922,WX8919,WX8920);
	or 	XG14361 	(WX8929,WX8926,WX8927);
	or 	XG14362 	(WX8936,WX8933,WX8934);
	or 	XG14363 	(WX8943,WX8940,WX8941);
	or 	XG14364 	(WX8950,WX8947,WX8948);
	or 	XG14365 	(WX8957,WX8954,WX8955);
	or 	XG14366 	(WX8964,WX8961,WX8962);
	or 	XG14367 	(WX8971,WX8968,WX8969);
	or 	XG14368 	(WX8978,WX8975,WX8976);
	or 	XG14369 	(WX8985,WX8982,WX8983);
	or 	XG14370 	(WX10061,WX10058,WX10059);
	or 	XG14371 	(WX10068,WX10065,WX10066);
	or 	XG14372 	(WX10075,WX10072,WX10073);
	or 	XG14373 	(WX10082,WX10079,WX10080);
	or 	XG14374 	(WX10089,WX10086,WX10087);
	or 	XG14375 	(WX10096,WX10093,WX10094);
	or 	XG14376 	(WX10103,WX10100,WX10101);
	or 	XG14377 	(WX10110,WX10107,WX10108);
	or 	XG14378 	(WX10117,WX10114,WX10115);
	or 	XG14379 	(WX10124,WX10121,WX10122);
	or 	XG14380 	(WX10131,WX10128,WX10129);
	or 	XG14381 	(WX10138,WX10135,WX10136);
	or 	XG14382 	(WX10145,WX10142,WX10143);
	or 	XG14383 	(WX10152,WX10149,WX10150);
	or 	XG14384 	(WX10159,WX10156,WX10157);
	or 	XG14385 	(WX10166,WX10163,WX10164);
	or 	XG14386 	(WX10173,WX10170,WX10171);
	or 	XG14387 	(WX10180,WX10177,WX10178);
	or 	XG14388 	(WX10187,WX10184,WX10185);
	or 	XG14389 	(WX10194,WX10191,WX10192);
	or 	XG14390 	(WX10201,WX10198,WX10199);
	or 	XG14391 	(WX10208,WX10205,WX10206);
	or 	XG14392 	(WX10215,WX10212,WX10213);
	or 	XG14393 	(WX10222,WX10219,WX10220);
	or 	XG14394 	(WX10229,WX10226,WX10227);
	or 	XG14395 	(WX10236,WX10233,WX10234);
	or 	XG14396 	(WX10243,WX10240,WX10241);
	or 	XG14397 	(WX10250,WX10247,WX10248);
	or 	XG14398 	(WX10257,WX10254,WX10255);
	or 	XG14399 	(WX10264,WX10261,WX10262);
	or 	XG14400 	(WX10271,WX10268,WX10269);
	or 	XG14401 	(WX10278,WX10275,WX10276);
	or 	XG14402 	(WX11354,WX11351,WX11352);
	or 	XG14403 	(WX11361,WX11358,WX11359);
	or 	XG14404 	(WX11368,WX11365,WX11366);
	or 	XG14405 	(WX11375,WX11372,WX11373);
	or 	XG14406 	(WX11382,WX11379,WX11380);
	or 	XG14407 	(WX11389,WX11386,WX11387);
	or 	XG14408 	(WX11396,WX11393,WX11394);
	or 	XG14409 	(WX11403,WX11400,WX11401);
	or 	XG14410 	(WX11410,WX11407,WX11408);
	or 	XG14411 	(WX11417,WX11414,WX11415);
	or 	XG14412 	(WX11424,WX11421,WX11422);
	or 	XG14413 	(WX11431,WX11428,WX11429);
	or 	XG14414 	(WX11438,WX11435,WX11436);
	or 	XG14415 	(WX11445,WX11442,WX11443);
	or 	XG14416 	(WX11452,WX11449,WX11450);
	or 	XG14417 	(WX11459,WX11456,WX11457);
	or 	XG14418 	(WX11466,WX11463,WX11464);
	or 	XG14419 	(WX11473,WX11470,WX11471);
	or 	XG14420 	(WX11480,WX11477,WX11478);
	or 	XG14421 	(WX11487,WX11484,WX11485);
	or 	XG14422 	(WX11494,WX11491,WX11492);
	or 	XG14423 	(WX11501,WX11498,WX11499);
	or 	XG14424 	(WX11508,WX11505,WX11506);
	or 	XG14425 	(WX11515,WX11512,WX11513);
	or 	XG14426 	(WX11522,WX11519,WX11520);
	or 	XG14427 	(WX11529,WX11526,WX11527);
	or 	XG14428 	(WX11536,WX11533,WX11534);
	or 	XG14429 	(WX11543,WX11540,WX11541);
	or 	XG14430 	(WX11550,WX11547,WX11548);
	or 	XG14431 	(WX11557,WX11554,WX11555);
	or 	XG14432 	(WX11564,WX11561,WX11562);
	or 	XG14433 	(WX11571,WX11568,WX11569);
	not 	XG14434 	(WX11572,WX11571);
	not 	XG14435 	(WX11565,WX11564);
	not 	XG14436 	(WX11558,WX11557);
	not 	XG14437 	(WX11551,WX11550);
	not 	XG14438 	(WX11544,WX11543);
	not 	XG14439 	(WX11537,WX11536);
	not 	XG14440 	(WX11530,WX11529);
	not 	XG14441 	(WX11523,WX11522);
	not 	XG14442 	(WX11516,WX11515);
	not 	XG14443 	(WX11509,WX11508);
	not 	XG14444 	(WX11502,WX11501);
	not 	XG14445 	(WX11495,WX11494);
	not 	XG14446 	(WX11488,WX11487);
	not 	XG14447 	(WX11481,WX11480);
	not 	XG14448 	(WX11474,WX11473);
	not 	XG14449 	(WX11467,WX11466);
	not 	XG14450 	(WX11460,WX11459);
	not 	XG14451 	(WX11453,WX11452);
	not 	XG14452 	(WX11446,WX11445);
	not 	XG14453 	(WX11439,WX11438);
	not 	XG14454 	(WX11432,WX11431);
	not 	XG14455 	(WX11425,WX11424);
	not 	XG14456 	(WX11418,WX11417);
	not 	XG14457 	(WX11411,WX11410);
	not 	XG14458 	(WX11404,WX11403);
	not 	XG14459 	(WX11397,WX11396);
	not 	XG14460 	(WX11390,WX11389);
	not 	XG14461 	(WX11383,WX11382);
	not 	XG14462 	(WX11376,WX11375);
	not 	XG14463 	(WX11369,WX11368);
	not 	XG14464 	(WX11362,WX11361);
	not 	XG14465 	(WX11355,WX11354);
	not 	XG14466 	(WX10279,WX10278);
	not 	XG14467 	(WX10272,WX10271);
	not 	XG14468 	(WX10265,WX10264);
	not 	XG14469 	(WX10258,WX10257);
	not 	XG14470 	(WX10251,WX10250);
	not 	XG14471 	(WX10244,WX10243);
	not 	XG14472 	(WX10237,WX10236);
	not 	XG14473 	(WX10230,WX10229);
	not 	XG14474 	(WX10223,WX10222);
	not 	XG14475 	(WX10216,WX10215);
	not 	XG14476 	(WX10209,WX10208);
	not 	XG14477 	(WX10202,WX10201);
	not 	XG14478 	(WX10195,WX10194);
	not 	XG14479 	(WX10188,WX10187);
	not 	XG14480 	(WX10181,WX10180);
	not 	XG14481 	(WX10174,WX10173);
	not 	XG14482 	(WX10167,WX10166);
	not 	XG14483 	(WX10160,WX10159);
	not 	XG14484 	(WX10153,WX10152);
	not 	XG14485 	(WX10146,WX10145);
	not 	XG14486 	(WX10139,WX10138);
	not 	XG14487 	(WX10132,WX10131);
	not 	XG14488 	(WX10125,WX10124);
	not 	XG14489 	(WX10118,WX10117);
	not 	XG14490 	(WX10111,WX10110);
	not 	XG14491 	(WX10104,WX10103);
	not 	XG14492 	(WX10097,WX10096);
	not 	XG14493 	(WX10090,WX10089);
	not 	XG14494 	(WX10083,WX10082);
	not 	XG14495 	(WX10076,WX10075);
	not 	XG14496 	(WX10069,WX10068);
	not 	XG14497 	(WX10062,WX10061);
	not 	XG14498 	(WX8986,WX8985);
	not 	XG14499 	(WX8979,WX8978);
	not 	XG14500 	(WX8972,WX8971);
	not 	XG14501 	(WX8965,WX8964);
	not 	XG14502 	(WX8958,WX8957);
	not 	XG14503 	(WX8951,WX8950);
	not 	XG14504 	(WX8944,WX8943);
	not 	XG14505 	(WX8937,WX8936);
	not 	XG14506 	(WX8930,WX8929);
	not 	XG14507 	(WX8923,WX8922);
	not 	XG14508 	(WX8916,WX8915);
	not 	XG14509 	(WX8909,WX8908);
	not 	XG14510 	(WX8902,WX8901);
	not 	XG14511 	(WX8895,WX8894);
	not 	XG14512 	(WX8888,WX8887);
	not 	XG14513 	(WX8881,WX8880);
	not 	XG14514 	(WX8874,WX8873);
	not 	XG14515 	(WX8867,WX8866);
	not 	XG14516 	(WX8860,WX8859);
	not 	XG14517 	(WX8853,WX8852);
	not 	XG14518 	(WX8846,WX8845);
	not 	XG14519 	(WX8839,WX8838);
	not 	XG14520 	(WX8832,WX8831);
	not 	XG14521 	(WX8825,WX8824);
	not 	XG14522 	(WX8818,WX8817);
	not 	XG14523 	(WX8811,WX8810);
	not 	XG14524 	(WX8804,WX8803);
	not 	XG14525 	(WX8797,WX8796);
	not 	XG14526 	(WX8790,WX8789);
	not 	XG14527 	(WX8783,WX8782);
	not 	XG14528 	(WX8776,WX8775);
	not 	XG14529 	(WX8769,WX8768);
	not 	XG14530 	(WX7693,WX7692);
	not 	XG14531 	(WX7686,WX7685);
	not 	XG14532 	(WX7679,WX7678);
	not 	XG14533 	(WX7672,WX7671);
	not 	XG14534 	(WX7665,WX7664);
	not 	XG14535 	(WX7658,WX7657);
	not 	XG14536 	(WX7651,WX7650);
	not 	XG14537 	(WX7644,WX7643);
	not 	XG14538 	(WX7637,WX7636);
	not 	XG14539 	(WX7630,WX7629);
	not 	XG14540 	(WX7623,WX7622);
	not 	XG14541 	(WX7616,WX7615);
	not 	XG14542 	(WX7609,WX7608);
	not 	XG14543 	(WX7602,WX7601);
	not 	XG14544 	(WX7595,WX7594);
	not 	XG14545 	(WX7588,WX7587);
	not 	XG14546 	(WX7581,WX7580);
	not 	XG14547 	(WX7574,WX7573);
	not 	XG14548 	(WX7567,WX7566);
	not 	XG14549 	(WX7560,WX7559);
	not 	XG14550 	(WX7553,WX7552);
	not 	XG14551 	(WX7546,WX7545);
	not 	XG14552 	(WX7539,WX7538);
	not 	XG14553 	(WX7532,WX7531);
	not 	XG14554 	(WX7525,WX7524);
	not 	XG14555 	(WX7518,WX7517);
	not 	XG14556 	(WX7511,WX7510);
	not 	XG14557 	(WX7504,WX7503);
	not 	XG14558 	(WX7497,WX7496);
	not 	XG14559 	(WX7490,WX7489);
	not 	XG14560 	(WX7483,WX7482);
	not 	XG14561 	(WX7476,WX7475);
	not 	XG14562 	(WX6400,WX6399);
	not 	XG14563 	(WX6393,WX6392);
	not 	XG14564 	(WX6386,WX6385);
	not 	XG14565 	(WX6379,WX6378);
	not 	XG14566 	(WX6372,WX6371);
	not 	XG14567 	(WX6365,WX6364);
	not 	XG14568 	(WX6358,WX6357);
	not 	XG14569 	(WX6351,WX6350);
	not 	XG14570 	(WX6344,WX6343);
	not 	XG14571 	(WX6337,WX6336);
	not 	XG14572 	(WX6330,WX6329);
	not 	XG14573 	(WX6323,WX6322);
	not 	XG14574 	(WX6316,WX6315);
	not 	XG14575 	(WX6309,WX6308);
	not 	XG14576 	(WX6302,WX6301);
	not 	XG14577 	(WX6295,WX6294);
	not 	XG14578 	(WX6288,WX6287);
	not 	XG14579 	(WX6281,WX6280);
	not 	XG14580 	(WX6274,WX6273);
	not 	XG14581 	(WX6267,WX6266);
	not 	XG14582 	(WX6260,WX6259);
	not 	XG14583 	(WX6253,WX6252);
	not 	XG14584 	(WX6246,WX6245);
	not 	XG14585 	(WX6239,WX6238);
	not 	XG14586 	(WX6232,WX6231);
	not 	XG14587 	(WX6225,WX6224);
	not 	XG14588 	(WX6218,WX6217);
	not 	XG14589 	(WX6211,WX6210);
	not 	XG14590 	(WX6204,WX6203);
	not 	XG14591 	(WX6197,WX6196);
	not 	XG14592 	(WX6190,WX6189);
	not 	XG14593 	(WX6183,WX6182);
	not 	XG14594 	(WX5107,WX5106);
	not 	XG14595 	(WX5100,WX5099);
	not 	XG14596 	(WX5093,WX5092);
	not 	XG14597 	(WX5086,WX5085);
	not 	XG14598 	(WX5079,WX5078);
	not 	XG14599 	(WX5072,WX5071);
	not 	XG14600 	(WX5065,WX5064);
	not 	XG14601 	(WX5058,WX5057);
	not 	XG14602 	(WX5051,WX5050);
	not 	XG14603 	(WX5044,WX5043);
	not 	XG14604 	(WX5037,WX5036);
	not 	XG14605 	(WX5030,WX5029);
	not 	XG14606 	(WX5023,WX5022);
	not 	XG14607 	(WX5016,WX5015);
	not 	XG14608 	(WX5009,WX5008);
	not 	XG14609 	(WX5002,WX5001);
	not 	XG14610 	(WX4995,WX4994);
	not 	XG14611 	(WX4988,WX4987);
	not 	XG14612 	(WX4981,WX4980);
	not 	XG14613 	(WX4974,WX4973);
	not 	XG14614 	(WX4967,WX4966);
	not 	XG14615 	(WX4960,WX4959);
	not 	XG14616 	(WX4953,WX4952);
	not 	XG14617 	(WX4946,WX4945);
	not 	XG14618 	(WX4939,WX4938);
	not 	XG14619 	(WX4932,WX4931);
	not 	XG14620 	(WX4925,WX4924);
	not 	XG14621 	(WX4918,WX4917);
	not 	XG14622 	(WX4911,WX4910);
	not 	XG14623 	(WX4904,WX4903);
	not 	XG14624 	(WX4897,WX4896);
	not 	XG14625 	(WX4890,WX4889);
	not 	XG14626 	(WX3814,WX3813);
	not 	XG14627 	(WX3807,WX3806);
	not 	XG14628 	(WX3800,WX3799);
	not 	XG14629 	(WX3793,WX3792);
	not 	XG14630 	(WX3786,WX3785);
	not 	XG14631 	(WX3779,WX3778);
	not 	XG14632 	(WX3772,WX3771);
	not 	XG14633 	(WX3765,WX3764);
	not 	XG14634 	(WX3758,WX3757);
	not 	XG14635 	(WX3751,WX3750);
	not 	XG14636 	(WX3744,WX3743);
	not 	XG14637 	(WX3737,WX3736);
	not 	XG14638 	(WX3730,WX3729);
	not 	XG14639 	(WX3723,WX3722);
	not 	XG14640 	(WX3716,WX3715);
	not 	XG14641 	(WX3709,WX3708);
	not 	XG14642 	(WX3702,WX3701);
	not 	XG14643 	(WX3695,WX3694);
	not 	XG14644 	(WX3688,WX3687);
	not 	XG14645 	(WX3681,WX3680);
	not 	XG14646 	(WX3674,WX3673);
	not 	XG14647 	(WX3667,WX3666);
	not 	XG14648 	(WX3660,WX3659);
	not 	XG14649 	(WX3653,WX3652);
	not 	XG14650 	(WX3646,WX3645);
	not 	XG14651 	(WX3639,WX3638);
	not 	XG14652 	(WX3632,WX3631);
	not 	XG14653 	(WX3625,WX3624);
	not 	XG14654 	(WX3618,WX3617);
	not 	XG14655 	(WX3611,WX3610);
	not 	XG14656 	(WX3604,WX3603);
	not 	XG14657 	(WX3597,WX3596);
	not 	XG14658 	(WX2521,WX2520);
	not 	XG14659 	(WX2514,WX2513);
	not 	XG14660 	(WX2507,WX2506);
	not 	XG14661 	(WX2500,WX2499);
	not 	XG14662 	(WX2493,WX2492);
	not 	XG14663 	(WX2486,WX2485);
	not 	XG14664 	(WX2479,WX2478);
	not 	XG14665 	(WX2472,WX2471);
	not 	XG14666 	(WX2465,WX2464);
	not 	XG14667 	(WX2458,WX2457);
	not 	XG14668 	(WX2451,WX2450);
	not 	XG14669 	(WX2444,WX2443);
	not 	XG14670 	(WX2437,WX2436);
	not 	XG14671 	(WX2430,WX2429);
	not 	XG14672 	(WX2423,WX2422);
	not 	XG14673 	(WX2416,WX2415);
	not 	XG14674 	(WX2409,WX2408);
	not 	XG14675 	(WX2402,WX2401);
	not 	XG14676 	(WX2395,WX2394);
	not 	XG14677 	(WX2388,WX2387);
	not 	XG14678 	(WX2381,WX2380);
	not 	XG14679 	(WX2374,WX2373);
	not 	XG14680 	(WX2367,WX2366);
	not 	XG14681 	(WX2360,WX2359);
	not 	XG14682 	(WX2353,WX2352);
	not 	XG14683 	(WX2346,WX2345);
	not 	XG14684 	(WX2339,WX2338);
	not 	XG14685 	(WX2332,WX2331);
	not 	XG14686 	(WX2325,WX2324);
	not 	XG14687 	(WX2318,WX2317);
	not 	XG14688 	(WX2311,WX2310);
	not 	XG14689 	(WX2304,WX2303);
	not 	XG14690 	(WX1228,WX1227);
	not 	XG14691 	(WX1221,WX1220);
	not 	XG14692 	(WX1214,WX1213);
	not 	XG14693 	(WX1207,WX1206);
	not 	XG14694 	(WX1200,WX1199);
	not 	XG14695 	(WX1193,WX1192);
	not 	XG14696 	(WX1186,WX1185);
	not 	XG14697 	(WX1179,WX1178);
	not 	XG14698 	(WX1172,WX1171);
	not 	XG14699 	(WX1165,WX1164);
	not 	XG14700 	(WX1158,WX1157);
	not 	XG14701 	(WX1151,WX1150);
	not 	XG14702 	(WX1144,WX1143);
	not 	XG14703 	(WX1137,WX1136);
	not 	XG14704 	(WX1130,WX1129);
	not 	XG14705 	(WX1123,WX1122);
	not 	XG14706 	(WX1116,WX1115);
	not 	XG14707 	(WX1109,WX1108);
	not 	XG14708 	(WX1102,WX1101);
	not 	XG14709 	(WX1095,WX1094);
	not 	XG14710 	(WX1088,WX1087);
	not 	XG14711 	(WX1081,WX1080);
	not 	XG14712 	(WX1074,WX1073);
	not 	XG14713 	(WX1067,WX1066);
	not 	XG14714 	(WX1060,WX1059);
	not 	XG14715 	(WX1053,WX1052);
	not 	XG14716 	(WX1046,WX1045);
	not 	XG14717 	(WX1039,WX1038);
	not 	XG14718 	(WX1032,WX1031);
	not 	XG14719 	(WX1025,WX1024);
	not 	XG14720 	(WX1018,WX1017);
	not 	XG14721 	(WX1011,WX1010);
	not 	XG14722 	(DATA_9_31,WX1011);
	not 	XG14723 	(DATA_9_30,WX1018);
	not 	XG14724 	(DATA_9_29,WX1025);
	not 	XG14725 	(DATA_9_28,WX1032);
	not 	XG14726 	(DATA_9_27,WX1039);
	not 	XG14727 	(DATA_9_26,WX1046);
	not 	XG14728 	(DATA_9_25,WX1053);
	not 	XG14729 	(DATA_9_24,WX1060);
	not 	XG14730 	(DATA_9_23,WX1067);
	not 	XG14731 	(DATA_9_22,WX1074);
	not 	XG14732 	(DATA_9_21,WX1081);
	not 	XG14733 	(DATA_9_20,WX1088);
	not 	XG14734 	(DATA_9_19,WX1095);
	not 	XG14735 	(DATA_9_18,WX1102);
	not 	XG14736 	(DATA_9_17,WX1109);
	not 	XG14737 	(DATA_9_16,WX1116);
	not 	XG14738 	(DATA_9_15,WX1123);
	not 	XG14739 	(DATA_9_14,WX1130);
	not 	XG14740 	(DATA_9_13,WX1137);
	not 	XG14741 	(DATA_9_12,WX1144);
	not 	XG14742 	(DATA_9_11,WX1151);
	not 	XG14743 	(DATA_9_10,WX1158);
	not 	XG14744 	(DATA_9_9,WX1165);
	not 	XG14745 	(DATA_9_8,WX1172);
	not 	XG14746 	(DATA_9_7,WX1179);
	not 	XG14747 	(DATA_9_6,WX1186);
	not 	XG14748 	(DATA_9_5,WX1193);
	not 	XG14749 	(DATA_9_4,WX1200);
	not 	XG14750 	(DATA_9_3,WX1207);
	not 	XG14751 	(DATA_9_2,WX1214);
	not 	XG14752 	(DATA_9_1,WX1221);
	not 	XG14753 	(DATA_9_0,WX1228);
	not 	XG14754 	(WX2305,WX2304);
	not 	XG14755 	(WX2312,WX2311);
	not 	XG14756 	(WX2319,WX2318);
	not 	XG14757 	(WX2326,WX2325);
	not 	XG14758 	(WX2333,WX2332);
	not 	XG14759 	(WX2340,WX2339);
	not 	XG14760 	(WX2347,WX2346);
	not 	XG14761 	(WX2354,WX2353);
	not 	XG14762 	(WX2361,WX2360);
	not 	XG14763 	(WX2368,WX2367);
	not 	XG14764 	(WX2375,WX2374);
	not 	XG14765 	(WX2382,WX2381);
	not 	XG14766 	(WX2389,WX2388);
	not 	XG14767 	(WX2396,WX2395);
	not 	XG14768 	(WX2403,WX2402);
	not 	XG14769 	(WX2410,WX2409);
	not 	XG14770 	(WX2417,WX2416);
	not 	XG14771 	(WX2424,WX2423);
	not 	XG14772 	(WX2431,WX2430);
	not 	XG14773 	(WX2438,WX2437);
	not 	XG14774 	(WX2445,WX2444);
	not 	XG14775 	(WX2452,WX2451);
	not 	XG14776 	(WX2459,WX2458);
	not 	XG14777 	(WX2466,WX2465);
	not 	XG14778 	(WX2473,WX2472);
	not 	XG14779 	(WX2480,WX2479);
	not 	XG14780 	(WX2487,WX2486);
	not 	XG14781 	(WX2494,WX2493);
	not 	XG14782 	(WX2501,WX2500);
	not 	XG14783 	(WX2508,WX2507);
	not 	XG14784 	(WX2515,WX2514);
	not 	XG14785 	(WX2522,WX2521);
	not 	XG14786 	(WX3598,WX3597);
	not 	XG14787 	(WX3605,WX3604);
	not 	XG14788 	(WX3612,WX3611);
	not 	XG14789 	(WX3619,WX3618);
	not 	XG14790 	(WX3626,WX3625);
	not 	XG14791 	(WX3633,WX3632);
	not 	XG14792 	(WX3640,WX3639);
	not 	XG14793 	(WX3647,WX3646);
	not 	XG14794 	(WX3654,WX3653);
	not 	XG14795 	(WX3661,WX3660);
	not 	XG14796 	(WX3668,WX3667);
	not 	XG14797 	(WX3675,WX3674);
	not 	XG14798 	(WX3682,WX3681);
	not 	XG14799 	(WX3689,WX3688);
	not 	XG14800 	(WX3696,WX3695);
	not 	XG14801 	(WX3703,WX3702);
	not 	XG14802 	(WX3710,WX3709);
	not 	XG14803 	(WX3717,WX3716);
	not 	XG14804 	(WX3724,WX3723);
	not 	XG14805 	(WX3731,WX3730);
	not 	XG14806 	(WX3738,WX3737);
	not 	XG14807 	(WX3745,WX3744);
	not 	XG14808 	(WX3752,WX3751);
	not 	XG14809 	(WX3759,WX3758);
	not 	XG14810 	(WX3766,WX3765);
	not 	XG14811 	(WX3773,WX3772);
	not 	XG14812 	(WX3780,WX3779);
	not 	XG14813 	(WX3787,WX3786);
	not 	XG14814 	(WX3794,WX3793);
	not 	XG14815 	(WX3801,WX3800);
	not 	XG14816 	(WX3808,WX3807);
	not 	XG14817 	(WX3815,WX3814);
	not 	XG14818 	(WX4891,WX4890);
	not 	XG14819 	(WX4898,WX4897);
	not 	XG14820 	(WX4905,WX4904);
	not 	XG14821 	(WX4912,WX4911);
	not 	XG14822 	(WX4919,WX4918);
	not 	XG14823 	(WX4926,WX4925);
	not 	XG14824 	(WX4933,WX4932);
	not 	XG14825 	(WX4940,WX4939);
	not 	XG14826 	(WX4947,WX4946);
	not 	XG14827 	(WX4954,WX4953);
	not 	XG14828 	(WX4961,WX4960);
	not 	XG14829 	(WX4968,WX4967);
	not 	XG14830 	(WX4975,WX4974);
	not 	XG14831 	(WX4982,WX4981);
	not 	XG14832 	(WX4989,WX4988);
	not 	XG14833 	(WX4996,WX4995);
	not 	XG14834 	(WX5003,WX5002);
	not 	XG14835 	(WX5010,WX5009);
	not 	XG14836 	(WX5017,WX5016);
	not 	XG14837 	(WX5024,WX5023);
	not 	XG14838 	(WX5031,WX5030);
	not 	XG14839 	(WX5038,WX5037);
	not 	XG14840 	(WX5045,WX5044);
	not 	XG14841 	(WX5052,WX5051);
	not 	XG14842 	(WX5059,WX5058);
	not 	XG14843 	(WX5066,WX5065);
	not 	XG14844 	(WX5073,WX5072);
	not 	XG14845 	(WX5080,WX5079);
	not 	XG14846 	(WX5087,WX5086);
	not 	XG14847 	(WX5094,WX5093);
	not 	XG14848 	(WX5101,WX5100);
	not 	XG14849 	(WX5108,WX5107);
	not 	XG14850 	(WX6184,WX6183);
	not 	XG14851 	(WX6191,WX6190);
	not 	XG14852 	(WX6198,WX6197);
	not 	XG14853 	(WX6205,WX6204);
	not 	XG14854 	(WX6212,WX6211);
	not 	XG14855 	(WX6219,WX6218);
	not 	XG14856 	(WX6226,WX6225);
	not 	XG14857 	(WX6233,WX6232);
	not 	XG14858 	(WX6240,WX6239);
	not 	XG14859 	(WX6247,WX6246);
	not 	XG14860 	(WX6254,WX6253);
	not 	XG14861 	(WX6261,WX6260);
	not 	XG14862 	(WX6268,WX6267);
	not 	XG14863 	(WX6275,WX6274);
	not 	XG14864 	(WX6282,WX6281);
	not 	XG14865 	(WX6289,WX6288);
	not 	XG14866 	(WX6296,WX6295);
	not 	XG14867 	(WX6303,WX6302);
	not 	XG14868 	(WX6310,WX6309);
	not 	XG14869 	(WX6317,WX6316);
	not 	XG14870 	(WX6324,WX6323);
	not 	XG14871 	(WX6331,WX6330);
	not 	XG14872 	(WX6338,WX6337);
	not 	XG14873 	(WX6345,WX6344);
	not 	XG14874 	(WX6352,WX6351);
	not 	XG14875 	(WX6359,WX6358);
	not 	XG14876 	(WX6366,WX6365);
	not 	XG14877 	(WX6373,WX6372);
	not 	XG14878 	(WX6380,WX6379);
	not 	XG14879 	(WX6387,WX6386);
	not 	XG14880 	(WX6394,WX6393);
	not 	XG14881 	(WX6401,WX6400);
	not 	XG14882 	(WX7477,WX7476);
	not 	XG14883 	(WX7484,WX7483);
	not 	XG14884 	(WX7491,WX7490);
	not 	XG14885 	(WX7498,WX7497);
	not 	XG14886 	(WX7505,WX7504);
	not 	XG14887 	(WX7512,WX7511);
	not 	XG14888 	(WX7519,WX7518);
	not 	XG14889 	(WX7526,WX7525);
	not 	XG14890 	(WX7533,WX7532);
	not 	XG14891 	(WX7540,WX7539);
	not 	XG14892 	(WX7547,WX7546);
	not 	XG14893 	(WX7554,WX7553);
	not 	XG14894 	(WX7561,WX7560);
	not 	XG14895 	(WX7568,WX7567);
	not 	XG14896 	(WX7575,WX7574);
	not 	XG14897 	(WX7582,WX7581);
	not 	XG14898 	(WX7589,WX7588);
	not 	XG14899 	(WX7596,WX7595);
	not 	XG14900 	(WX7603,WX7602);
	not 	XG14901 	(WX7610,WX7609);
	not 	XG14902 	(WX7617,WX7616);
	not 	XG14903 	(WX7624,WX7623);
	not 	XG14904 	(WX7631,WX7630);
	not 	XG14905 	(WX7638,WX7637);
	not 	XG14906 	(WX7645,WX7644);
	not 	XG14907 	(WX7652,WX7651);
	not 	XG14908 	(WX7659,WX7658);
	not 	XG14909 	(WX7666,WX7665);
	not 	XG14910 	(WX7673,WX7672);
	not 	XG14911 	(WX7680,WX7679);
	not 	XG14912 	(WX7687,WX7686);
	not 	XG14913 	(WX7694,WX7693);
	not 	XG14914 	(WX8770,WX8769);
	not 	XG14915 	(WX8777,WX8776);
	not 	XG14916 	(WX8784,WX8783);
	not 	XG14917 	(WX8791,WX8790);
	not 	XG14918 	(WX8798,WX8797);
	not 	XG14919 	(WX8805,WX8804);
	not 	XG14920 	(WX8812,WX8811);
	not 	XG14921 	(WX8819,WX8818);
	not 	XG14922 	(WX8826,WX8825);
	not 	XG14923 	(WX8833,WX8832);
	not 	XG14924 	(WX8840,WX8839);
	not 	XG14925 	(WX8847,WX8846);
	not 	XG14926 	(WX8854,WX8853);
	not 	XG14927 	(WX8861,WX8860);
	not 	XG14928 	(WX8868,WX8867);
	not 	XG14929 	(WX8875,WX8874);
	not 	XG14930 	(WX8882,WX8881);
	not 	XG14931 	(WX8889,WX8888);
	not 	XG14932 	(WX8896,WX8895);
	not 	XG14933 	(WX8903,WX8902);
	not 	XG14934 	(WX8910,WX8909);
	not 	XG14935 	(WX8917,WX8916);
	not 	XG14936 	(WX8924,WX8923);
	not 	XG14937 	(WX8931,WX8930);
	not 	XG14938 	(WX8938,WX8937);
	not 	XG14939 	(WX8945,WX8944);
	not 	XG14940 	(WX8952,WX8951);
	not 	XG14941 	(WX8959,WX8958);
	not 	XG14942 	(WX8966,WX8965);
	not 	XG14943 	(WX8973,WX8972);
	not 	XG14944 	(WX8980,WX8979);
	not 	XG14945 	(WX8987,WX8986);
	not 	XG14946 	(WX10063,WX10062);
	not 	XG14947 	(WX10070,WX10069);
	not 	XG14948 	(WX10077,WX10076);
	not 	XG14949 	(WX10084,WX10083);
	not 	XG14950 	(WX10091,WX10090);
	not 	XG14951 	(WX10098,WX10097);
	not 	XG14952 	(WX10105,WX10104);
	not 	XG14953 	(WX10112,WX10111);
	not 	XG14954 	(WX10119,WX10118);
	not 	XG14955 	(WX10126,WX10125);
	not 	XG14956 	(WX10133,WX10132);
	not 	XG14957 	(WX10140,WX10139);
	not 	XG14958 	(WX10147,WX10146);
	not 	XG14959 	(WX10154,WX10153);
	not 	XG14960 	(WX10161,WX10160);
	not 	XG14961 	(WX10168,WX10167);
	not 	XG14962 	(WX10175,WX10174);
	not 	XG14963 	(WX10182,WX10181);
	not 	XG14964 	(WX10189,WX10188);
	not 	XG14965 	(WX10196,WX10195);
	not 	XG14966 	(WX10203,WX10202);
	not 	XG14967 	(WX10210,WX10209);
	not 	XG14968 	(WX10217,WX10216);
	not 	XG14969 	(WX10224,WX10223);
	not 	XG14970 	(WX10231,WX10230);
	not 	XG14971 	(WX10238,WX10237);
	not 	XG14972 	(WX10245,WX10244);
	not 	XG14973 	(WX10252,WX10251);
	not 	XG14974 	(WX10259,WX10258);
	not 	XG14975 	(WX10266,WX10265);
	not 	XG14976 	(WX10273,WX10272);
	not 	XG14977 	(WX10280,WX10279);
	not 	XG14978 	(WX11356,WX11355);
	not 	XG14979 	(WX11363,WX11362);
	not 	XG14980 	(WX11370,WX11369);
	not 	XG14981 	(WX11377,WX11376);
	not 	XG14982 	(WX11384,WX11383);
	not 	XG14983 	(WX11391,WX11390);
	not 	XG14984 	(WX11398,WX11397);
	not 	XG14985 	(WX11405,WX11404);
	not 	XG14986 	(WX11412,WX11411);
	not 	XG14987 	(WX11419,WX11418);
	not 	XG14988 	(WX11426,WX11425);
	not 	XG14989 	(WX11433,WX11432);
	not 	XG14990 	(WX11440,WX11439);
	not 	XG14991 	(WX11447,WX11446);
	not 	XG14992 	(WX11454,WX11453);
	not 	XG14993 	(WX11461,WX11460);
	not 	XG14994 	(WX11468,WX11467);
	not 	XG14995 	(WX11475,WX11474);
	not 	XG14996 	(WX11482,WX11481);
	not 	XG14997 	(WX11489,WX11488);
	not 	XG14998 	(WX11496,WX11495);
	not 	XG14999 	(WX11503,WX11502);
	not 	XG15000 	(WX11510,WX11509);
	not 	XG15001 	(WX11517,WX11516);
	not 	XG15002 	(WX11524,WX11523);
	not 	XG15003 	(WX11531,WX11530);
	not 	XG15004 	(WX11538,WX11537);
	not 	XG15005 	(WX11545,WX11544);
	not 	XG15006 	(WX11552,WX11551);
	not 	XG15007 	(WX11559,WX11558);
	not 	XG15008 	(WX11566,WX11565);
	not 	XG15009 	(WX11573,WX11572);
	and 	XG15010 	(WX10822,WX10823,WX11573);
	and 	XG15011 	(WX10808,WX10809,WX11566);
	and 	XG15012 	(WX10794,WX10795,WX11559);
	and 	XG15013 	(WX10780,WX10781,WX11552);
	and 	XG15014 	(WX10766,WX10767,WX11545);
	and 	XG15015 	(WX10752,WX10753,WX11538);
	and 	XG15016 	(WX10738,WX10739,WX11531);
	and 	XG15017 	(WX10724,WX10725,WX11524);
	and 	XG15018 	(WX10710,WX10711,WX11517);
	and 	XG15019 	(WX10696,WX10697,WX11510);
	and 	XG15020 	(WX10682,WX10683,WX11503);
	and 	XG15021 	(WX10668,WX10669,WX11496);
	and 	XG15022 	(WX10654,WX10655,WX11489);
	and 	XG15023 	(WX10640,WX10641,WX11482);
	and 	XG15024 	(WX10626,WX10627,WX11475);
	and 	XG15025 	(WX10612,WX10613,WX11468);
	and 	XG15026 	(WX10598,WX10599,WX11461);
	and 	XG15027 	(WX10584,WX10585,WX11454);
	and 	XG15028 	(WX10570,WX10571,WX11447);
	and 	XG15029 	(WX10556,WX10557,WX11440);
	and 	XG15030 	(WX10542,WX10543,WX11433);
	and 	XG15031 	(WX10528,WX10529,WX11426);
	and 	XG15032 	(WX10514,WX10515,WX11419);
	and 	XG15033 	(WX10500,WX10501,WX11412);
	and 	XG15034 	(WX10486,WX10487,WX11405);
	and 	XG15035 	(WX10472,WX10473,WX11398);
	and 	XG15036 	(WX10458,WX10459,WX11391);
	and 	XG15037 	(WX10444,WX10445,WX11384);
	and 	XG15038 	(WX10430,WX10431,WX11377);
	and 	XG15039 	(WX10416,WX10417,WX11370);
	and 	XG15040 	(WX10402,WX10403,WX11363);
	and 	XG15041 	(WX10388,WX10389,WX11356);
	and 	XG15042 	(WX9529,WX9530,WX10280);
	and 	XG15043 	(WX9515,WX9516,WX10273);
	and 	XG15044 	(WX9501,WX9502,WX10266);
	and 	XG15045 	(WX9487,WX9488,WX10259);
	and 	XG15046 	(WX9473,WX9474,WX10252);
	and 	XG15047 	(WX9459,WX9460,WX10245);
	and 	XG15048 	(WX9445,WX9446,WX10238);
	and 	XG15049 	(WX9431,WX9432,WX10231);
	and 	XG15050 	(WX9417,WX9418,WX10224);
	and 	XG15051 	(WX9403,WX9404,WX10217);
	and 	XG15052 	(WX9389,WX9390,WX10210);
	and 	XG15053 	(WX9375,WX9376,WX10203);
	and 	XG15054 	(WX9361,WX9362,WX10196);
	and 	XG15055 	(WX9347,WX9348,WX10189);
	and 	XG15056 	(WX9333,WX9334,WX10182);
	and 	XG15057 	(WX9319,WX9320,WX10175);
	and 	XG15058 	(WX9305,WX9306,WX10168);
	and 	XG15059 	(WX9291,WX9292,WX10161);
	and 	XG15060 	(WX9277,WX9278,WX10154);
	and 	XG15061 	(WX9263,WX9264,WX10147);
	and 	XG15062 	(WX9249,WX9250,WX10140);
	and 	XG15063 	(WX9235,WX9236,WX10133);
	and 	XG15064 	(WX9221,WX9222,WX10126);
	and 	XG15065 	(WX9207,WX9208,WX10119);
	and 	XG15066 	(WX9193,WX9194,WX10112);
	and 	XG15067 	(WX9179,WX9180,WX10105);
	and 	XG15068 	(WX9165,WX9166,WX10098);
	and 	XG15069 	(WX9151,WX9152,WX10091);
	and 	XG15070 	(WX9137,WX9138,WX10084);
	and 	XG15071 	(WX9123,WX9124,WX10077);
	and 	XG15072 	(WX9109,WX9110,WX10070);
	and 	XG15073 	(WX9095,WX9096,WX10063);
	and 	XG15074 	(WX8236,WX8237,WX8987);
	and 	XG15075 	(WX8222,WX8223,WX8980);
	and 	XG15076 	(WX8208,WX8209,WX8973);
	and 	XG15077 	(WX8194,WX8195,WX8966);
	and 	XG15078 	(WX8180,WX8181,WX8959);
	and 	XG15079 	(WX8166,WX8167,WX8952);
	and 	XG15080 	(WX8152,WX8153,WX8945);
	and 	XG15081 	(WX8138,WX8139,WX8938);
	and 	XG15082 	(WX8124,WX8125,WX8931);
	and 	XG15083 	(WX8110,WX8111,WX8924);
	and 	XG15084 	(WX8096,WX8097,WX8917);
	and 	XG15085 	(WX8082,WX8083,WX8910);
	and 	XG15086 	(WX8068,WX8069,WX8903);
	and 	XG15087 	(WX8054,WX8055,WX8896);
	and 	XG15088 	(WX8040,WX8041,WX8889);
	and 	XG15089 	(WX8026,WX8027,WX8882);
	and 	XG15090 	(WX8012,WX8013,WX8875);
	and 	XG15091 	(WX7998,WX7999,WX8868);
	and 	XG15092 	(WX7984,WX7985,WX8861);
	and 	XG15093 	(WX7970,WX7971,WX8854);
	and 	XG15094 	(WX7956,WX7957,WX8847);
	and 	XG15095 	(WX7942,WX7943,WX8840);
	and 	XG15096 	(WX7928,WX7929,WX8833);
	and 	XG15097 	(WX7914,WX7915,WX8826);
	and 	XG15098 	(WX7900,WX7901,WX8819);
	and 	XG15099 	(WX7886,WX7887,WX8812);
	and 	XG15100 	(WX7872,WX7873,WX8805);
	and 	XG15101 	(WX7858,WX7859,WX8798);
	and 	XG15102 	(WX7844,WX7845,WX8791);
	and 	XG15103 	(WX7830,WX7831,WX8784);
	and 	XG15104 	(WX7816,WX7817,WX8777);
	and 	XG15105 	(WX7802,WX7803,WX8770);
	and 	XG15106 	(WX6943,WX6944,WX7694);
	and 	XG15107 	(WX6929,WX6930,WX7687);
	and 	XG15108 	(WX6915,WX6916,WX7680);
	and 	XG15109 	(WX6901,WX6902,WX7673);
	and 	XG15110 	(WX6887,WX6888,WX7666);
	and 	XG15111 	(WX6873,WX6874,WX7659);
	and 	XG15112 	(WX6859,WX6860,WX7652);
	and 	XG15113 	(WX6845,WX6846,WX7645);
	and 	XG15114 	(WX6831,WX6832,WX7638);
	and 	XG15115 	(WX6817,WX6818,WX7631);
	and 	XG15116 	(WX6803,WX6804,WX7624);
	and 	XG15117 	(WX6789,WX6790,WX7617);
	and 	XG15118 	(WX6775,WX6776,WX7610);
	and 	XG15119 	(WX6761,WX6762,WX7603);
	and 	XG15120 	(WX6747,WX6748,WX7596);
	and 	XG15121 	(WX6733,WX6734,WX7589);
	and 	XG15122 	(WX6719,WX6720,WX7582);
	and 	XG15123 	(WX6705,WX6706,WX7575);
	and 	XG15124 	(WX6691,WX6692,WX7568);
	and 	XG15125 	(WX6677,WX6678,WX7561);
	and 	XG15126 	(WX6663,WX6664,WX7554);
	and 	XG15127 	(WX6649,WX6650,WX7547);
	and 	XG15128 	(WX6635,WX6636,WX7540);
	and 	XG15129 	(WX6621,WX6622,WX7533);
	and 	XG15130 	(WX6607,WX6608,WX7526);
	and 	XG15131 	(WX6593,WX6594,WX7519);
	and 	XG15132 	(WX6579,WX6580,WX7512);
	and 	XG15133 	(WX6565,WX6566,WX7505);
	and 	XG15134 	(WX6551,WX6552,WX7498);
	and 	XG15135 	(WX6537,WX6538,WX7491);
	and 	XG15136 	(WX6523,WX6524,WX7484);
	and 	XG15137 	(WX6509,WX6510,WX7477);
	and 	XG15138 	(WX5650,WX5651,WX6401);
	and 	XG15139 	(WX5636,WX5637,WX6394);
	and 	XG15140 	(WX5622,WX5623,WX6387);
	and 	XG15141 	(WX5608,WX5609,WX6380);
	and 	XG15142 	(WX5594,WX5595,WX6373);
	and 	XG15143 	(WX5580,WX5581,WX6366);
	and 	XG15144 	(WX5566,WX5567,WX6359);
	and 	XG15145 	(WX5552,WX5553,WX6352);
	and 	XG15146 	(WX5538,WX5539,WX6345);
	and 	XG15147 	(WX5524,WX5525,WX6338);
	and 	XG15148 	(WX5510,WX5511,WX6331);
	and 	XG15149 	(WX5496,WX5497,WX6324);
	and 	XG15150 	(WX5482,WX5483,WX6317);
	and 	XG15151 	(WX5468,WX5469,WX6310);
	and 	XG15152 	(WX5454,WX5455,WX6303);
	and 	XG15153 	(WX5440,WX5441,WX6296);
	and 	XG15154 	(WX5426,WX5427,WX6289);
	and 	XG15155 	(WX5412,WX5413,WX6282);
	and 	XG15156 	(WX5398,WX5399,WX6275);
	and 	XG15157 	(WX5384,WX5385,WX6268);
	and 	XG15158 	(WX5370,WX5371,WX6261);
	and 	XG15159 	(WX5356,WX5357,WX6254);
	and 	XG15160 	(WX5342,WX5343,WX6247);
	and 	XG15161 	(WX5328,WX5329,WX6240);
	and 	XG15162 	(WX5314,WX5315,WX6233);
	and 	XG15163 	(WX5300,WX5301,WX6226);
	and 	XG15164 	(WX5286,WX5287,WX6219);
	and 	XG15165 	(WX5272,WX5273,WX6212);
	and 	XG15166 	(WX5258,WX5259,WX6205);
	and 	XG15167 	(WX5244,WX5245,WX6198);
	and 	XG15168 	(WX5230,WX5231,WX6191);
	and 	XG15169 	(WX5216,WX5217,WX6184);
	and 	XG15170 	(WX4357,WX4358,WX5108);
	and 	XG15171 	(WX4343,WX4344,WX5101);
	and 	XG15172 	(WX4329,WX4330,WX5094);
	and 	XG15173 	(WX4315,WX4316,WX5087);
	and 	XG15174 	(WX4301,WX4302,WX5080);
	and 	XG15175 	(WX4287,WX4288,WX5073);
	and 	XG15176 	(WX4273,WX4274,WX5066);
	and 	XG15177 	(WX4259,WX4260,WX5059);
	and 	XG15178 	(WX4245,WX4246,WX5052);
	and 	XG15179 	(WX4231,WX4232,WX5045);
	and 	XG15180 	(WX4217,WX4218,WX5038);
	and 	XG15181 	(WX4203,WX4204,WX5031);
	and 	XG15182 	(WX4189,WX4190,WX5024);
	and 	XG15183 	(WX4175,WX4176,WX5017);
	and 	XG15184 	(WX4161,WX4162,WX5010);
	and 	XG15185 	(WX4147,WX4148,WX5003);
	and 	XG15186 	(WX4133,WX4134,WX4996);
	and 	XG15187 	(WX4119,WX4120,WX4989);
	and 	XG15188 	(WX4105,WX4106,WX4982);
	and 	XG15189 	(WX4091,WX4092,WX4975);
	and 	XG15190 	(WX4077,WX4078,WX4968);
	and 	XG15191 	(WX4063,WX4064,WX4961);
	and 	XG15192 	(WX4049,WX4050,WX4954);
	and 	XG15193 	(WX4035,WX4036,WX4947);
	and 	XG15194 	(WX4021,WX4022,WX4940);
	and 	XG15195 	(WX4007,WX4008,WX4933);
	and 	XG15196 	(WX3993,WX3994,WX4926);
	and 	XG15197 	(WX3979,WX3980,WX4919);
	and 	XG15198 	(WX3965,WX3966,WX4912);
	and 	XG15199 	(WX3951,WX3952,WX4905);
	and 	XG15200 	(WX3937,WX3938,WX4898);
	and 	XG15201 	(WX3923,WX3924,WX4891);
	and 	XG15202 	(WX3064,WX3065,WX3815);
	and 	XG15203 	(WX3050,WX3051,WX3808);
	and 	XG15204 	(WX3036,WX3037,WX3801);
	and 	XG15205 	(WX3022,WX3023,WX3794);
	and 	XG15206 	(WX3008,WX3009,WX3787);
	and 	XG15207 	(WX2994,WX2995,WX3780);
	and 	XG15208 	(WX2980,WX2981,WX3773);
	and 	XG15209 	(WX2966,WX2967,WX3766);
	and 	XG15210 	(WX2952,WX2953,WX3759);
	and 	XG15211 	(WX2938,WX2939,WX3752);
	and 	XG15212 	(WX2924,WX2925,WX3745);
	and 	XG15213 	(WX2910,WX2911,WX3738);
	and 	XG15214 	(WX2896,WX2897,WX3731);
	and 	XG15215 	(WX2882,WX2883,WX3724);
	and 	XG15216 	(WX2868,WX2869,WX3717);
	and 	XG15217 	(WX2854,WX2855,WX3710);
	and 	XG15218 	(WX2840,WX2841,WX3703);
	and 	XG15219 	(WX2826,WX2827,WX3696);
	and 	XG15220 	(WX2812,WX2813,WX3689);
	and 	XG15221 	(WX2798,WX2799,WX3682);
	and 	XG15222 	(WX2784,WX2785,WX3675);
	and 	XG15223 	(WX2770,WX2771,WX3668);
	and 	XG15224 	(WX2756,WX2757,WX3661);
	and 	XG15225 	(WX2742,WX2743,WX3654);
	and 	XG15226 	(WX2728,WX2729,WX3647);
	and 	XG15227 	(WX2714,WX2715,WX3640);
	and 	XG15228 	(WX2700,WX2701,WX3633);
	and 	XG15229 	(WX2686,WX2687,WX3626);
	and 	XG15230 	(WX2672,WX2673,WX3619);
	and 	XG15231 	(WX2658,WX2659,WX3612);
	and 	XG15232 	(WX2644,WX2645,WX3605);
	and 	XG15233 	(WX2630,WX2631,WX3598);
	and 	XG15234 	(WX1771,WX1772,WX2522);
	and 	XG15235 	(WX1757,WX1758,WX2515);
	and 	XG15236 	(WX1743,WX1744,WX2508);
	and 	XG15237 	(WX1729,WX1730,WX2501);
	and 	XG15238 	(WX1715,WX1716,WX2494);
	and 	XG15239 	(WX1701,WX1702,WX2487);
	and 	XG15240 	(WX1687,WX1688,WX2480);
	and 	XG15241 	(WX1673,WX1674,WX2473);
	and 	XG15242 	(WX1659,WX1660,WX2466);
	and 	XG15243 	(WX1645,WX1646,WX2459);
	and 	XG15244 	(WX1631,WX1632,WX2452);
	and 	XG15245 	(WX1617,WX1618,WX2445);
	and 	XG15246 	(WX1603,WX1604,WX2438);
	and 	XG15247 	(WX1589,WX1590,WX2431);
	and 	XG15248 	(WX1575,WX1576,WX2424);
	and 	XG15249 	(WX1561,WX1562,WX2417);
	and 	XG15250 	(WX1547,WX1548,WX2410);
	and 	XG15251 	(WX1533,WX1534,WX2403);
	and 	XG15252 	(WX1519,WX1520,WX2396);
	and 	XG15253 	(WX1505,WX1506,WX2389);
	and 	XG15254 	(WX1491,WX1492,WX2382);
	and 	XG15255 	(WX1477,WX1478,WX2375);
	and 	XG15256 	(WX1463,WX1464,WX2368);
	and 	XG15257 	(WX1449,WX1450,WX2361);
	and 	XG15258 	(WX1435,WX1436,WX2354);
	and 	XG15259 	(WX1421,WX1422,WX2347);
	and 	XG15260 	(WX1407,WX1408,WX2340);
	and 	XG15261 	(WX1393,WX1394,WX2333);
	and 	XG15262 	(WX1379,WX1380,WX2326);
	and 	XG15263 	(WX1365,WX1366,WX2319);
	and 	XG15264 	(WX1351,WX1352,WX2312);
	and 	XG15265 	(WX1337,WX1338,WX2305);
	and 	XG15266 	(WX478,WX479,DATA_9_0);
	and 	XG15267 	(WX464,WX465,DATA_9_1);
	and 	XG15268 	(WX450,WX451,DATA_9_2);
	and 	XG15269 	(WX436,WX437,DATA_9_3);
	and 	XG15270 	(WX422,WX423,DATA_9_4);
	and 	XG15271 	(WX408,WX409,DATA_9_5);
	and 	XG15272 	(WX394,WX395,DATA_9_6);
	and 	XG15273 	(WX380,WX381,DATA_9_7);
	and 	XG15274 	(WX366,WX367,DATA_9_8);
	and 	XG15275 	(WX352,WX353,DATA_9_9);
	and 	XG15276 	(WX338,WX339,DATA_9_10);
	and 	XG15277 	(WX324,WX325,DATA_9_11);
	and 	XG15278 	(WX310,WX311,DATA_9_12);
	and 	XG15279 	(WX296,WX297,DATA_9_13);
	and 	XG15280 	(WX282,WX283,DATA_9_14);
	and 	XG15281 	(WX268,WX269,DATA_9_15);
	and 	XG15282 	(WX254,WX255,DATA_9_16);
	and 	XG15283 	(WX240,WX241,DATA_9_17);
	and 	XG15284 	(WX226,WX227,DATA_9_18);
	and 	XG15285 	(WX212,WX213,DATA_9_19);
	and 	XG15286 	(WX198,WX199,DATA_9_20);
	and 	XG15287 	(WX184,WX185,DATA_9_21);
	and 	XG15288 	(WX170,WX171,DATA_9_22);
	and 	XG15289 	(WX156,WX157,DATA_9_23);
	and 	XG15290 	(WX142,WX143,DATA_9_24);
	and 	XG15291 	(WX128,WX129,DATA_9_25);
	and 	XG15292 	(WX114,WX115,DATA_9_26);
	and 	XG15293 	(WX100,WX101,DATA_9_27);
	and 	XG15294 	(WX86,WX87,DATA_9_28);
	and 	XG15295 	(WX72,WX73,DATA_9_29);
	and 	XG15296 	(WX58,WX59,DATA_9_30);
	and 	XG15297 	(WX44,WX45,DATA_9_31);
	and 	XG15298 	(WX40,WX41,WX2305);
	and 	XG15299 	(WX54,WX55,WX2312);
	and 	XG15300 	(WX68,WX69,WX2319);
	and 	XG15301 	(WX82,WX83,WX2326);
	and 	XG15302 	(WX96,WX97,WX2333);
	and 	XG15303 	(WX110,WX111,WX2340);
	and 	XG15304 	(WX124,WX125,WX2347);
	and 	XG15305 	(WX138,WX139,WX2354);
	and 	XG15306 	(WX152,WX153,WX2361);
	and 	XG15307 	(WX166,WX167,WX2368);
	and 	XG15308 	(WX180,WX181,WX2375);
	and 	XG15309 	(WX194,WX195,WX2382);
	and 	XG15310 	(WX208,WX209,WX2389);
	and 	XG15311 	(WX222,WX223,WX2396);
	and 	XG15312 	(WX236,WX237,WX2403);
	and 	XG15313 	(WX250,WX251,WX2410);
	and 	XG15314 	(WX264,WX265,WX2417);
	and 	XG15315 	(WX278,WX279,WX2424);
	and 	XG15316 	(WX292,WX293,WX2431);
	and 	XG15317 	(WX306,WX307,WX2438);
	and 	XG15318 	(WX320,WX321,WX2445);
	and 	XG15319 	(WX334,WX335,WX2452);
	and 	XG15320 	(WX348,WX349,WX2459);
	and 	XG15321 	(WX362,WX363,WX2466);
	and 	XG15322 	(WX376,WX377,WX2473);
	and 	XG15323 	(WX390,WX391,WX2480);
	and 	XG15324 	(WX404,WX405,WX2487);
	and 	XG15325 	(WX418,WX419,WX2494);
	and 	XG15326 	(WX432,WX433,WX2501);
	and 	XG15327 	(WX446,WX447,WX2508);
	and 	XG15328 	(WX460,WX461,WX2515);
	and 	XG15329 	(WX474,WX475,WX2522);
	and 	XG15330 	(WX1333,WX1334,WX3598);
	and 	XG15331 	(WX1347,WX1348,WX3605);
	and 	XG15332 	(WX1361,WX1362,WX3612);
	and 	XG15333 	(WX1375,WX1376,WX3619);
	and 	XG15334 	(WX1389,WX1390,WX3626);
	and 	XG15335 	(WX1403,WX1404,WX3633);
	and 	XG15336 	(WX1417,WX1418,WX3640);
	and 	XG15337 	(WX1431,WX1432,WX3647);
	and 	XG15338 	(WX1445,WX1446,WX3654);
	and 	XG15339 	(WX1459,WX1460,WX3661);
	and 	XG15340 	(WX1473,WX1474,WX3668);
	and 	XG15341 	(WX1487,WX1488,WX3675);
	and 	XG15342 	(WX1501,WX1502,WX3682);
	and 	XG15343 	(WX1515,WX1516,WX3689);
	and 	XG15344 	(WX1529,WX1530,WX3696);
	and 	XG15345 	(WX1543,WX1544,WX3703);
	and 	XG15346 	(WX1557,WX1558,WX3710);
	and 	XG15347 	(WX1571,WX1572,WX3717);
	and 	XG15348 	(WX1585,WX1586,WX3724);
	and 	XG15349 	(WX1599,WX1600,WX3731);
	and 	XG15350 	(WX1613,WX1614,WX3738);
	and 	XG15351 	(WX1627,WX1628,WX3745);
	and 	XG15352 	(WX1641,WX1642,WX3752);
	and 	XG15353 	(WX1655,WX1656,WX3759);
	and 	XG15354 	(WX1669,WX1670,WX3766);
	and 	XG15355 	(WX1683,WX1684,WX3773);
	and 	XG15356 	(WX1697,WX1698,WX3780);
	and 	XG15357 	(WX1711,WX1712,WX3787);
	and 	XG15358 	(WX1725,WX1726,WX3794);
	and 	XG15359 	(WX1739,WX1740,WX3801);
	and 	XG15360 	(WX1753,WX1754,WX3808);
	and 	XG15361 	(WX1767,WX1768,WX3815);
	and 	XG15362 	(WX2626,WX2627,WX4891);
	and 	XG15363 	(WX2640,WX2641,WX4898);
	and 	XG15364 	(WX2654,WX2655,WX4905);
	and 	XG15365 	(WX2668,WX2669,WX4912);
	and 	XG15366 	(WX2682,WX2683,WX4919);
	and 	XG15367 	(WX2696,WX2697,WX4926);
	and 	XG15368 	(WX2710,WX2711,WX4933);
	and 	XG15369 	(WX2724,WX2725,WX4940);
	and 	XG15370 	(WX2738,WX2739,WX4947);
	and 	XG15371 	(WX2752,WX2753,WX4954);
	and 	XG15372 	(WX2766,WX2767,WX4961);
	and 	XG15373 	(WX2780,WX2781,WX4968);
	and 	XG15374 	(WX2794,WX2795,WX4975);
	and 	XG15375 	(WX2808,WX2809,WX4982);
	and 	XG15376 	(WX2822,WX2823,WX4989);
	and 	XG15377 	(WX2836,WX2837,WX4996);
	and 	XG15378 	(WX2850,WX2851,WX5003);
	and 	XG15379 	(WX2864,WX2865,WX5010);
	and 	XG15380 	(WX2878,WX2879,WX5017);
	and 	XG15381 	(WX2892,WX2893,WX5024);
	and 	XG15382 	(WX2906,WX2907,WX5031);
	and 	XG15383 	(WX2920,WX2921,WX5038);
	and 	XG15384 	(WX2934,WX2935,WX5045);
	and 	XG15385 	(WX2948,WX2949,WX5052);
	and 	XG15386 	(WX2962,WX2963,WX5059);
	and 	XG15387 	(WX2976,WX2977,WX5066);
	and 	XG15388 	(WX2990,WX2991,WX5073);
	and 	XG15389 	(WX3004,WX3005,WX5080);
	and 	XG15390 	(WX3018,WX3019,WX5087);
	and 	XG15391 	(WX3032,WX3033,WX5094);
	and 	XG15392 	(WX3046,WX3047,WX5101);
	and 	XG15393 	(WX3060,WX3061,WX5108);
	and 	XG15394 	(WX3919,WX3920,WX6184);
	and 	XG15395 	(WX3933,WX3934,WX6191);
	and 	XG15396 	(WX3947,WX3948,WX6198);
	and 	XG15397 	(WX3961,WX3962,WX6205);
	and 	XG15398 	(WX3975,WX3976,WX6212);
	and 	XG15399 	(WX3989,WX3990,WX6219);
	and 	XG15400 	(WX4003,WX4004,WX6226);
	and 	XG15401 	(WX4017,WX4018,WX6233);
	and 	XG15402 	(WX4031,WX4032,WX6240);
	and 	XG15403 	(WX4045,WX4046,WX6247);
	and 	XG15404 	(WX4059,WX4060,WX6254);
	and 	XG15405 	(WX4073,WX4074,WX6261);
	and 	XG15406 	(WX4087,WX4088,WX6268);
	and 	XG15407 	(WX4101,WX4102,WX6275);
	and 	XG15408 	(WX4115,WX4116,WX6282);
	and 	XG15409 	(WX4129,WX4130,WX6289);
	and 	XG15410 	(WX4143,WX4144,WX6296);
	and 	XG15411 	(WX4157,WX4158,WX6303);
	and 	XG15412 	(WX4171,WX4172,WX6310);
	and 	XG15413 	(WX4185,WX4186,WX6317);
	and 	XG15414 	(WX4199,WX4200,WX6324);
	and 	XG15415 	(WX4213,WX4214,WX6331);
	and 	XG15416 	(WX4227,WX4228,WX6338);
	and 	XG15417 	(WX4241,WX4242,WX6345);
	and 	XG15418 	(WX4255,WX4256,WX6352);
	and 	XG15419 	(WX4269,WX4270,WX6359);
	and 	XG15420 	(WX4283,WX4284,WX6366);
	and 	XG15421 	(WX4297,WX4298,WX6373);
	and 	XG15422 	(WX4311,WX4312,WX6380);
	and 	XG15423 	(WX4325,WX4326,WX6387);
	and 	XG15424 	(WX4339,WX4340,WX6394);
	and 	XG15425 	(WX4353,WX4354,WX6401);
	and 	XG15426 	(WX5212,WX5213,WX7477);
	and 	XG15427 	(WX5226,WX5227,WX7484);
	and 	XG15428 	(WX5240,WX5241,WX7491);
	and 	XG15429 	(WX5254,WX5255,WX7498);
	and 	XG15430 	(WX5268,WX5269,WX7505);
	and 	XG15431 	(WX5282,WX5283,WX7512);
	and 	XG15432 	(WX5296,WX5297,WX7519);
	and 	XG15433 	(WX5310,WX5311,WX7526);
	and 	XG15434 	(WX5324,WX5325,WX7533);
	and 	XG15435 	(WX5338,WX5339,WX7540);
	and 	XG15436 	(WX5352,WX5353,WX7547);
	and 	XG15437 	(WX5366,WX5367,WX7554);
	and 	XG15438 	(WX5380,WX5381,WX7561);
	and 	XG15439 	(WX5394,WX5395,WX7568);
	and 	XG15440 	(WX5408,WX5409,WX7575);
	and 	XG15441 	(WX5422,WX5423,WX7582);
	and 	XG15442 	(WX5436,WX5437,WX7589);
	and 	XG15443 	(WX5450,WX5451,WX7596);
	and 	XG15444 	(WX5464,WX5465,WX7603);
	and 	XG15445 	(WX5478,WX5479,WX7610);
	and 	XG15446 	(WX5492,WX5493,WX7617);
	and 	XG15447 	(WX5506,WX5507,WX7624);
	and 	XG15448 	(WX5520,WX5521,WX7631);
	and 	XG15449 	(WX5534,WX5535,WX7638);
	and 	XG15450 	(WX5548,WX5549,WX7645);
	and 	XG15451 	(WX5562,WX5563,WX7652);
	and 	XG15452 	(WX5576,WX5577,WX7659);
	and 	XG15453 	(WX5590,WX5591,WX7666);
	and 	XG15454 	(WX5604,WX5605,WX7673);
	and 	XG15455 	(WX5618,WX5619,WX7680);
	and 	XG15456 	(WX5632,WX5633,WX7687);
	and 	XG15457 	(WX5646,WX5647,WX7694);
	and 	XG15458 	(WX6505,WX6506,WX8770);
	and 	XG15459 	(WX6519,WX6520,WX8777);
	and 	XG15460 	(WX6533,WX6534,WX8784);
	and 	XG15461 	(WX6547,WX6548,WX8791);
	and 	XG15462 	(WX6561,WX6562,WX8798);
	and 	XG15463 	(WX6575,WX6576,WX8805);
	and 	XG15464 	(WX6589,WX6590,WX8812);
	and 	XG15465 	(WX6603,WX6604,WX8819);
	and 	XG15466 	(WX6617,WX6618,WX8826);
	and 	XG15467 	(WX6631,WX6632,WX8833);
	and 	XG15468 	(WX6645,WX6646,WX8840);
	and 	XG15469 	(WX6659,WX6660,WX8847);
	and 	XG15470 	(WX6673,WX6674,WX8854);
	and 	XG15471 	(WX6687,WX6688,WX8861);
	and 	XG15472 	(WX6701,WX6702,WX8868);
	and 	XG15473 	(WX6715,WX6716,WX8875);
	and 	XG15474 	(WX6729,WX6730,WX8882);
	and 	XG15475 	(WX6743,WX6744,WX8889);
	and 	XG15476 	(WX6757,WX6758,WX8896);
	and 	XG15477 	(WX6771,WX6772,WX8903);
	and 	XG15478 	(WX6785,WX6786,WX8910);
	and 	XG15479 	(WX6799,WX6800,WX8917);
	and 	XG15480 	(WX6813,WX6814,WX8924);
	and 	XG15481 	(WX6827,WX6828,WX8931);
	and 	XG15482 	(WX6841,WX6842,WX8938);
	and 	XG15483 	(WX6855,WX6856,WX8945);
	and 	XG15484 	(WX6869,WX6870,WX8952);
	and 	XG15485 	(WX6883,WX6884,WX8959);
	and 	XG15486 	(WX6897,WX6898,WX8966);
	and 	XG15487 	(WX6911,WX6912,WX8973);
	and 	XG15488 	(WX6925,WX6926,WX8980);
	and 	XG15489 	(WX6939,WX6940,WX8987);
	and 	XG15490 	(WX7798,WX7799,WX10063);
	and 	XG15491 	(WX7812,WX7813,WX10070);
	and 	XG15492 	(WX7826,WX7827,WX10077);
	and 	XG15493 	(WX7840,WX7841,WX10084);
	and 	XG15494 	(WX7854,WX7855,WX10091);
	and 	XG15495 	(WX7868,WX7869,WX10098);
	and 	XG15496 	(WX7882,WX7883,WX10105);
	and 	XG15497 	(WX7896,WX7897,WX10112);
	and 	XG15498 	(WX7910,WX7911,WX10119);
	and 	XG15499 	(WX7924,WX7925,WX10126);
	and 	XG15500 	(WX7938,WX7939,WX10133);
	and 	XG15501 	(WX7952,WX7953,WX10140);
	and 	XG15502 	(WX7966,WX7967,WX10147);
	and 	XG15503 	(WX7980,WX7981,WX10154);
	and 	XG15504 	(WX7994,WX7995,WX10161);
	and 	XG15505 	(WX8008,WX8009,WX10168);
	and 	XG15506 	(WX8022,WX8023,WX10175);
	and 	XG15507 	(WX8036,WX8037,WX10182);
	and 	XG15508 	(WX8050,WX8051,WX10189);
	and 	XG15509 	(WX8064,WX8065,WX10196);
	and 	XG15510 	(WX8078,WX8079,WX10203);
	and 	XG15511 	(WX8092,WX8093,WX10210);
	and 	XG15512 	(WX8106,WX8107,WX10217);
	and 	XG15513 	(WX8120,WX8121,WX10224);
	and 	XG15514 	(WX8134,WX8135,WX10231);
	and 	XG15515 	(WX8148,WX8149,WX10238);
	and 	XG15516 	(WX8162,WX8163,WX10245);
	and 	XG15517 	(WX8176,WX8177,WX10252);
	and 	XG15518 	(WX8190,WX8191,WX10259);
	and 	XG15519 	(WX8204,WX8205,WX10266);
	and 	XG15520 	(WX8218,WX8219,WX10273);
	and 	XG15521 	(WX8232,WX8233,WX10280);
	and 	XG15522 	(WX9091,WX9092,WX11356);
	and 	XG15523 	(WX9105,WX9106,WX11363);
	and 	XG15524 	(WX9119,WX9120,WX11370);
	and 	XG15525 	(WX9133,WX9134,WX11377);
	and 	XG15526 	(WX9147,WX9148,WX11384);
	and 	XG15527 	(WX9161,WX9162,WX11391);
	and 	XG15528 	(WX9175,WX9176,WX11398);
	and 	XG15529 	(WX9189,WX9190,WX11405);
	and 	XG15530 	(WX9203,WX9204,WX11412);
	and 	XG15531 	(WX9217,WX9218,WX11419);
	and 	XG15532 	(WX9231,WX9232,WX11426);
	and 	XG15533 	(WX9245,WX9246,WX11433);
	and 	XG15534 	(WX9259,WX9260,WX11440);
	and 	XG15535 	(WX9273,WX9274,WX11447);
	and 	XG15536 	(WX9287,WX9288,WX11454);
	and 	XG15537 	(WX9301,WX9302,WX11461);
	and 	XG15538 	(WX9315,WX9316,WX11468);
	and 	XG15539 	(WX9329,WX9330,WX11475);
	and 	XG15540 	(WX9343,WX9344,WX11482);
	and 	XG15541 	(WX9357,WX9358,WX11489);
	and 	XG15542 	(WX9371,WX9372,WX11496);
	and 	XG15543 	(WX9385,WX9386,WX11503);
	and 	XG15544 	(WX9399,WX9400,WX11510);
	and 	XG15545 	(WX9413,WX9414,WX11517);
	and 	XG15546 	(WX9427,WX9428,WX11524);
	and 	XG15547 	(WX9441,WX9442,WX11531);
	and 	XG15548 	(WX9455,WX9456,WX11538);
	and 	XG15549 	(WX9469,WX9470,WX11545);
	and 	XG15550 	(WX9483,WX9484,WX11552);
	and 	XG15551 	(WX9497,WX9498,WX11559);
	and 	XG15552 	(WX9511,WX9512,WX11566);
	and 	XG15553 	(WX9525,WX9526,WX11573);
	or 	XG15554 	(WX10824,WX10821,WX10822);
	or 	XG15555 	(WX10810,WX10807,WX10808);
	or 	XG15556 	(WX10796,WX10793,WX10794);
	or 	XG15557 	(WX10782,WX10779,WX10780);
	or 	XG15558 	(WX10768,WX10765,WX10766);
	or 	XG15559 	(WX10754,WX10751,WX10752);
	or 	XG15560 	(WX10740,WX10737,WX10738);
	or 	XG15561 	(WX10726,WX10723,WX10724);
	or 	XG15562 	(WX10712,WX10709,WX10710);
	or 	XG15563 	(WX10698,WX10695,WX10696);
	or 	XG15564 	(WX10684,WX10681,WX10682);
	or 	XG15565 	(WX10670,WX10667,WX10668);
	or 	XG15566 	(WX10656,WX10653,WX10654);
	or 	XG15567 	(WX10642,WX10639,WX10640);
	or 	XG15568 	(WX10628,WX10625,WX10626);
	or 	XG15569 	(WX10614,WX10611,WX10612);
	or 	XG15570 	(WX10600,WX10597,WX10598);
	or 	XG15571 	(WX10586,WX10583,WX10584);
	or 	XG15572 	(WX10572,WX10569,WX10570);
	or 	XG15573 	(WX10558,WX10555,WX10556);
	or 	XG15574 	(WX10544,WX10541,WX10542);
	or 	XG15575 	(WX10530,WX10527,WX10528);
	or 	XG15576 	(WX10516,WX10513,WX10514);
	or 	XG15577 	(WX10502,WX10499,WX10500);
	or 	XG15578 	(WX10488,WX10485,WX10486);
	or 	XG15579 	(WX10474,WX10471,WX10472);
	or 	XG15580 	(WX10460,WX10457,WX10458);
	or 	XG15581 	(WX10446,WX10443,WX10444);
	or 	XG15582 	(WX10432,WX10429,WX10430);
	or 	XG15583 	(WX10418,WX10415,WX10416);
	or 	XG15584 	(WX10404,WX10401,WX10402);
	or 	XG15585 	(WX10390,WX10387,WX10388);
	or 	XG15586 	(WX9531,WX9528,WX9529);
	or 	XG15587 	(WX9517,WX9514,WX9515);
	or 	XG15588 	(WX9503,WX9500,WX9501);
	or 	XG15589 	(WX9489,WX9486,WX9487);
	or 	XG15590 	(WX9475,WX9472,WX9473);
	or 	XG15591 	(WX9461,WX9458,WX9459);
	or 	XG15592 	(WX9447,WX9444,WX9445);
	or 	XG15593 	(WX9433,WX9430,WX9431);
	or 	XG15594 	(WX9419,WX9416,WX9417);
	or 	XG15595 	(WX9405,WX9402,WX9403);
	or 	XG15596 	(WX9391,WX9388,WX9389);
	or 	XG15597 	(WX9377,WX9374,WX9375);
	or 	XG15598 	(WX9363,WX9360,WX9361);
	or 	XG15599 	(WX9349,WX9346,WX9347);
	or 	XG15600 	(WX9335,WX9332,WX9333);
	or 	XG15601 	(WX9321,WX9318,WX9319);
	or 	XG15602 	(WX9307,WX9304,WX9305);
	or 	XG15603 	(WX9293,WX9290,WX9291);
	or 	XG15604 	(WX9279,WX9276,WX9277);
	or 	XG15605 	(WX9265,WX9262,WX9263);
	or 	XG15606 	(WX9251,WX9248,WX9249);
	or 	XG15607 	(WX9237,WX9234,WX9235);
	or 	XG15608 	(WX9223,WX9220,WX9221);
	or 	XG15609 	(WX9209,WX9206,WX9207);
	or 	XG15610 	(WX9195,WX9192,WX9193);
	or 	XG15611 	(WX9181,WX9178,WX9179);
	or 	XG15612 	(WX9167,WX9164,WX9165);
	or 	XG15613 	(WX9153,WX9150,WX9151);
	or 	XG15614 	(WX9139,WX9136,WX9137);
	or 	XG15615 	(WX9125,WX9122,WX9123);
	or 	XG15616 	(WX9111,WX9108,WX9109);
	or 	XG15617 	(WX9097,WX9094,WX9095);
	or 	XG15618 	(WX8238,WX8235,WX8236);
	or 	XG15619 	(WX8224,WX8221,WX8222);
	or 	XG15620 	(WX8210,WX8207,WX8208);
	or 	XG15621 	(WX8196,WX8193,WX8194);
	or 	XG15622 	(WX8182,WX8179,WX8180);
	or 	XG15623 	(WX8168,WX8165,WX8166);
	or 	XG15624 	(WX8154,WX8151,WX8152);
	or 	XG15625 	(WX8140,WX8137,WX8138);
	or 	XG15626 	(WX8126,WX8123,WX8124);
	or 	XG15627 	(WX8112,WX8109,WX8110);
	or 	XG15628 	(WX8098,WX8095,WX8096);
	or 	XG15629 	(WX8084,WX8081,WX8082);
	or 	XG15630 	(WX8070,WX8067,WX8068);
	or 	XG15631 	(WX8056,WX8053,WX8054);
	or 	XG15632 	(WX8042,WX8039,WX8040);
	or 	XG15633 	(WX8028,WX8025,WX8026);
	or 	XG15634 	(WX8014,WX8011,WX8012);
	or 	XG15635 	(WX8000,WX7997,WX7998);
	or 	XG15636 	(WX7986,WX7983,WX7984);
	or 	XG15637 	(WX7972,WX7969,WX7970);
	or 	XG15638 	(WX7958,WX7955,WX7956);
	or 	XG15639 	(WX7944,WX7941,WX7942);
	or 	XG15640 	(WX7930,WX7927,WX7928);
	or 	XG15641 	(WX7916,WX7913,WX7914);
	or 	XG15642 	(WX7902,WX7899,WX7900);
	or 	XG15643 	(WX7888,WX7885,WX7886);
	or 	XG15644 	(WX7874,WX7871,WX7872);
	or 	XG15645 	(WX7860,WX7857,WX7858);
	or 	XG15646 	(WX7846,WX7843,WX7844);
	or 	XG15647 	(WX7832,WX7829,WX7830);
	or 	XG15648 	(WX7818,WX7815,WX7816);
	or 	XG15649 	(WX7804,WX7801,WX7802);
	or 	XG15650 	(WX6945,WX6942,WX6943);
	or 	XG15651 	(WX6931,WX6928,WX6929);
	or 	XG15652 	(WX6917,WX6914,WX6915);
	or 	XG15653 	(WX6903,WX6900,WX6901);
	or 	XG15654 	(WX6889,WX6886,WX6887);
	or 	XG15655 	(WX6875,WX6872,WX6873);
	or 	XG15656 	(WX6861,WX6858,WX6859);
	or 	XG15657 	(WX6847,WX6844,WX6845);
	or 	XG15658 	(WX6833,WX6830,WX6831);
	or 	XG15659 	(WX6819,WX6816,WX6817);
	or 	XG15660 	(WX6805,WX6802,WX6803);
	or 	XG15661 	(WX6791,WX6788,WX6789);
	or 	XG15662 	(WX6777,WX6774,WX6775);
	or 	XG15663 	(WX6763,WX6760,WX6761);
	or 	XG15664 	(WX6749,WX6746,WX6747);
	or 	XG15665 	(WX6735,WX6732,WX6733);
	or 	XG15666 	(WX6721,WX6718,WX6719);
	or 	XG15667 	(WX6707,WX6704,WX6705);
	or 	XG15668 	(WX6693,WX6690,WX6691);
	or 	XG15669 	(WX6679,WX6676,WX6677);
	or 	XG15670 	(WX6665,WX6662,WX6663);
	or 	XG15671 	(WX6651,WX6648,WX6649);
	or 	XG15672 	(WX6637,WX6634,WX6635);
	or 	XG15673 	(WX6623,WX6620,WX6621);
	or 	XG15674 	(WX6609,WX6606,WX6607);
	or 	XG15675 	(WX6595,WX6592,WX6593);
	or 	XG15676 	(WX6581,WX6578,WX6579);
	or 	XG15677 	(WX6567,WX6564,WX6565);
	or 	XG15678 	(WX6553,WX6550,WX6551);
	or 	XG15679 	(WX6539,WX6536,WX6537);
	or 	XG15680 	(WX6525,WX6522,WX6523);
	or 	XG15681 	(WX6511,WX6508,WX6509);
	or 	XG15682 	(WX5652,WX5649,WX5650);
	or 	XG15683 	(WX5638,WX5635,WX5636);
	or 	XG15684 	(WX5624,WX5621,WX5622);
	or 	XG15685 	(WX5610,WX5607,WX5608);
	or 	XG15686 	(WX5596,WX5593,WX5594);
	or 	XG15687 	(WX5582,WX5579,WX5580);
	or 	XG15688 	(WX5568,WX5565,WX5566);
	or 	XG15689 	(WX5554,WX5551,WX5552);
	or 	XG15690 	(WX5540,WX5537,WX5538);
	or 	XG15691 	(WX5526,WX5523,WX5524);
	or 	XG15692 	(WX5512,WX5509,WX5510);
	or 	XG15693 	(WX5498,WX5495,WX5496);
	or 	XG15694 	(WX5484,WX5481,WX5482);
	or 	XG15695 	(WX5470,WX5467,WX5468);
	or 	XG15696 	(WX5456,WX5453,WX5454);
	or 	XG15697 	(WX5442,WX5439,WX5440);
	or 	XG15698 	(WX5428,WX5425,WX5426);
	or 	XG15699 	(WX5414,WX5411,WX5412);
	or 	XG15700 	(WX5400,WX5397,WX5398);
	or 	XG15701 	(WX5386,WX5383,WX5384);
	or 	XG15702 	(WX5372,WX5369,WX5370);
	or 	XG15703 	(WX5358,WX5355,WX5356);
	or 	XG15704 	(WX5344,WX5341,WX5342);
	or 	XG15705 	(WX5330,WX5327,WX5328);
	or 	XG15706 	(WX5316,WX5313,WX5314);
	or 	XG15707 	(WX5302,WX5299,WX5300);
	or 	XG15708 	(WX5288,WX5285,WX5286);
	or 	XG15709 	(WX5274,WX5271,WX5272);
	or 	XG15710 	(WX5260,WX5257,WX5258);
	or 	XG15711 	(WX5246,WX5243,WX5244);
	or 	XG15712 	(WX5232,WX5229,WX5230);
	or 	XG15713 	(WX5218,WX5215,WX5216);
	or 	XG15714 	(WX4359,WX4356,WX4357);
	or 	XG15715 	(WX4345,WX4342,WX4343);
	or 	XG15716 	(WX4331,WX4328,WX4329);
	or 	XG15717 	(WX4317,WX4314,WX4315);
	or 	XG15718 	(WX4303,WX4300,WX4301);
	or 	XG15719 	(WX4289,WX4286,WX4287);
	or 	XG15720 	(WX4275,WX4272,WX4273);
	or 	XG15721 	(WX4261,WX4258,WX4259);
	or 	XG15722 	(WX4247,WX4244,WX4245);
	or 	XG15723 	(WX4233,WX4230,WX4231);
	or 	XG15724 	(WX4219,WX4216,WX4217);
	or 	XG15725 	(WX4205,WX4202,WX4203);
	or 	XG15726 	(WX4191,WX4188,WX4189);
	or 	XG15727 	(WX4177,WX4174,WX4175);
	or 	XG15728 	(WX4163,WX4160,WX4161);
	or 	XG15729 	(WX4149,WX4146,WX4147);
	or 	XG15730 	(WX4135,WX4132,WX4133);
	or 	XG15731 	(WX4121,WX4118,WX4119);
	or 	XG15732 	(WX4107,WX4104,WX4105);
	or 	XG15733 	(WX4093,WX4090,WX4091);
	or 	XG15734 	(WX4079,WX4076,WX4077);
	or 	XG15735 	(WX4065,WX4062,WX4063);
	or 	XG15736 	(WX4051,WX4048,WX4049);
	or 	XG15737 	(WX4037,WX4034,WX4035);
	or 	XG15738 	(WX4023,WX4020,WX4021);
	or 	XG15739 	(WX4009,WX4006,WX4007);
	or 	XG15740 	(WX3995,WX3992,WX3993);
	or 	XG15741 	(WX3981,WX3978,WX3979);
	or 	XG15742 	(WX3967,WX3964,WX3965);
	or 	XG15743 	(WX3953,WX3950,WX3951);
	or 	XG15744 	(WX3939,WX3936,WX3937);
	or 	XG15745 	(WX3925,WX3922,WX3923);
	or 	XG15746 	(WX3066,WX3063,WX3064);
	or 	XG15747 	(WX3052,WX3049,WX3050);
	or 	XG15748 	(WX3038,WX3035,WX3036);
	or 	XG15749 	(WX3024,WX3021,WX3022);
	or 	XG15750 	(WX3010,WX3007,WX3008);
	or 	XG15751 	(WX2996,WX2993,WX2994);
	or 	XG15752 	(WX2982,WX2979,WX2980);
	or 	XG15753 	(WX2968,WX2965,WX2966);
	or 	XG15754 	(WX2954,WX2951,WX2952);
	or 	XG15755 	(WX2940,WX2937,WX2938);
	or 	XG15756 	(WX2926,WX2923,WX2924);
	or 	XG15757 	(WX2912,WX2909,WX2910);
	or 	XG15758 	(WX2898,WX2895,WX2896);
	or 	XG15759 	(WX2884,WX2881,WX2882);
	or 	XG15760 	(WX2870,WX2867,WX2868);
	or 	XG15761 	(WX2856,WX2853,WX2854);
	or 	XG15762 	(WX2842,WX2839,WX2840);
	or 	XG15763 	(WX2828,WX2825,WX2826);
	or 	XG15764 	(WX2814,WX2811,WX2812);
	or 	XG15765 	(WX2800,WX2797,WX2798);
	or 	XG15766 	(WX2786,WX2783,WX2784);
	or 	XG15767 	(WX2772,WX2769,WX2770);
	or 	XG15768 	(WX2758,WX2755,WX2756);
	or 	XG15769 	(WX2744,WX2741,WX2742);
	or 	XG15770 	(WX2730,WX2727,WX2728);
	or 	XG15771 	(WX2716,WX2713,WX2714);
	or 	XG15772 	(WX2702,WX2699,WX2700);
	or 	XG15773 	(WX2688,WX2685,WX2686);
	or 	XG15774 	(WX2674,WX2671,WX2672);
	or 	XG15775 	(WX2660,WX2657,WX2658);
	or 	XG15776 	(WX2646,WX2643,WX2644);
	or 	XG15777 	(WX2632,WX2629,WX2630);
	or 	XG15778 	(WX1773,WX1770,WX1771);
	or 	XG15779 	(WX1759,WX1756,WX1757);
	or 	XG15780 	(WX1745,WX1742,WX1743);
	or 	XG15781 	(WX1731,WX1728,WX1729);
	or 	XG15782 	(WX1717,WX1714,WX1715);
	or 	XG15783 	(WX1703,WX1700,WX1701);
	or 	XG15784 	(WX1689,WX1686,WX1687);
	or 	XG15785 	(WX1675,WX1672,WX1673);
	or 	XG15786 	(WX1661,WX1658,WX1659);
	or 	XG15787 	(WX1647,WX1644,WX1645);
	or 	XG15788 	(WX1633,WX1630,WX1631);
	or 	XG15789 	(WX1619,WX1616,WX1617);
	or 	XG15790 	(WX1605,WX1602,WX1603);
	or 	XG15791 	(WX1591,WX1588,WX1589);
	or 	XG15792 	(WX1577,WX1574,WX1575);
	or 	XG15793 	(WX1563,WX1560,WX1561);
	or 	XG15794 	(WX1549,WX1546,WX1547);
	or 	XG15795 	(WX1535,WX1532,WX1533);
	or 	XG15796 	(WX1521,WX1518,WX1519);
	or 	XG15797 	(WX1507,WX1504,WX1505);
	or 	XG15798 	(WX1493,WX1490,WX1491);
	or 	XG15799 	(WX1479,WX1476,WX1477);
	or 	XG15800 	(WX1465,WX1462,WX1463);
	or 	XG15801 	(WX1451,WX1448,WX1449);
	or 	XG15802 	(WX1437,WX1434,WX1435);
	or 	XG15803 	(WX1423,WX1420,WX1421);
	or 	XG15804 	(WX1409,WX1406,WX1407);
	or 	XG15805 	(WX1395,WX1392,WX1393);
	or 	XG15806 	(WX1381,WX1378,WX1379);
	or 	XG15807 	(WX1367,WX1364,WX1365);
	or 	XG15808 	(WX1353,WX1350,WX1351);
	or 	XG15809 	(WX1339,WX1336,WX1337);
	or 	XG15810 	(WX480,WX477,WX478);
	or 	XG15811 	(WX466,WX463,WX464);
	or 	XG15812 	(WX452,WX449,WX450);
	or 	XG15813 	(WX438,WX435,WX436);
	or 	XG15814 	(WX424,WX421,WX422);
	or 	XG15815 	(WX410,WX407,WX408);
	or 	XG15816 	(WX396,WX393,WX394);
	or 	XG15817 	(WX382,WX379,WX380);
	or 	XG15818 	(WX368,WX365,WX366);
	or 	XG15819 	(WX354,WX351,WX352);
	or 	XG15820 	(WX340,WX337,WX338);
	or 	XG15821 	(WX326,WX323,WX324);
	or 	XG15822 	(WX312,WX309,WX310);
	or 	XG15823 	(WX298,WX295,WX296);
	or 	XG15824 	(WX284,WX281,WX282);
	or 	XG15825 	(WX270,WX267,WX268);
	or 	XG15826 	(WX256,WX253,WX254);
	or 	XG15827 	(WX242,WX239,WX240);
	or 	XG15828 	(WX228,WX225,WX226);
	or 	XG15829 	(WX214,WX211,WX212);
	or 	XG15830 	(WX200,WX197,WX198);
	or 	XG15831 	(WX186,WX183,WX184);
	or 	XG15832 	(WX172,WX169,WX170);
	or 	XG15833 	(WX158,WX155,WX156);
	or 	XG15834 	(WX144,WX141,WX142);
	or 	XG15835 	(WX130,WX127,WX128);
	or 	XG15836 	(WX116,WX113,WX114);
	or 	XG15837 	(WX102,WX99,WX100);
	or 	XG15838 	(WX88,WX85,WX86);
	or 	XG15839 	(WX74,WX71,WX72);
	or 	XG15840 	(WX60,WX57,WX58);
	or 	XG15841 	(WX46,WX43,WX44);
	or 	XG15842 	(WX9093,WX9090,WX9091);
	or 	XG15843 	(WX9107,WX9104,WX9105);
	or 	XG15844 	(WX9121,WX9118,WX9119);
	or 	XG15845 	(WX9135,WX9132,WX9133);
	or 	XG15846 	(WX9149,WX9146,WX9147);
	or 	XG15847 	(WX9163,WX9160,WX9161);
	or 	XG15848 	(WX9177,WX9174,WX9175);
	or 	XG15849 	(WX9191,WX9188,WX9189);
	or 	XG15850 	(WX9205,WX9202,WX9203);
	or 	XG15851 	(WX9219,WX9216,WX9217);
	or 	XG15852 	(WX9233,WX9230,WX9231);
	or 	XG15853 	(WX9247,WX9244,WX9245);
	or 	XG15854 	(WX9261,WX9258,WX9259);
	or 	XG15855 	(WX9275,WX9272,WX9273);
	or 	XG15856 	(WX9289,WX9286,WX9287);
	or 	XG15857 	(WX9303,WX9300,WX9301);
	or 	XG15858 	(WX9317,WX9314,WX9315);
	or 	XG15859 	(WX9331,WX9328,WX9329);
	or 	XG15860 	(WX9345,WX9342,WX9343);
	or 	XG15861 	(WX9359,WX9356,WX9357);
	or 	XG15862 	(WX9373,WX9370,WX9371);
	or 	XG15863 	(WX9387,WX9384,WX9385);
	or 	XG15864 	(WX9401,WX9398,WX9399);
	or 	XG15865 	(WX9415,WX9412,WX9413);
	or 	XG15866 	(WX9429,WX9426,WX9427);
	or 	XG15867 	(WX9443,WX9440,WX9441);
	or 	XG15868 	(WX9457,WX9454,WX9455);
	or 	XG15869 	(WX9471,WX9468,WX9469);
	or 	XG15870 	(WX9485,WX9482,WX9483);
	or 	XG15871 	(WX9499,WX9496,WX9497);
	or 	XG15872 	(WX9513,WX9510,WX9511);
	or 	XG15873 	(WX9527,WX9524,WX9525);
	or 	XG15874 	(WX7800,WX7797,WX7798);
	or 	XG15875 	(WX7814,WX7811,WX7812);
	or 	XG15876 	(WX7828,WX7825,WX7826);
	or 	XG15877 	(WX7842,WX7839,WX7840);
	or 	XG15878 	(WX7856,WX7853,WX7854);
	or 	XG15879 	(WX7870,WX7867,WX7868);
	or 	XG15880 	(WX7884,WX7881,WX7882);
	or 	XG15881 	(WX7898,WX7895,WX7896);
	or 	XG15882 	(WX7912,WX7909,WX7910);
	or 	XG15883 	(WX7926,WX7923,WX7924);
	or 	XG15884 	(WX7940,WX7937,WX7938);
	or 	XG15885 	(WX7954,WX7951,WX7952);
	or 	XG15886 	(WX7968,WX7965,WX7966);
	or 	XG15887 	(WX7982,WX7979,WX7980);
	or 	XG15888 	(WX7996,WX7993,WX7994);
	or 	XG15889 	(WX8010,WX8007,WX8008);
	or 	XG15890 	(WX8024,WX8021,WX8022);
	or 	XG15891 	(WX8038,WX8035,WX8036);
	or 	XG15892 	(WX8052,WX8049,WX8050);
	or 	XG15893 	(WX8066,WX8063,WX8064);
	or 	XG15894 	(WX8080,WX8077,WX8078);
	or 	XG15895 	(WX8094,WX8091,WX8092);
	or 	XG15896 	(WX8108,WX8105,WX8106);
	or 	XG15897 	(WX8122,WX8119,WX8120);
	or 	XG15898 	(WX8136,WX8133,WX8134);
	or 	XG15899 	(WX8150,WX8147,WX8148);
	or 	XG15900 	(WX8164,WX8161,WX8162);
	or 	XG15901 	(WX8178,WX8175,WX8176);
	or 	XG15902 	(WX8192,WX8189,WX8190);
	or 	XG15903 	(WX8206,WX8203,WX8204);
	or 	XG15904 	(WX8220,WX8217,WX8218);
	or 	XG15905 	(WX8234,WX8231,WX8232);
	or 	XG15906 	(WX6507,WX6504,WX6505);
	or 	XG15907 	(WX6521,WX6518,WX6519);
	or 	XG15908 	(WX6535,WX6532,WX6533);
	or 	XG15909 	(WX6549,WX6546,WX6547);
	or 	XG15910 	(WX6563,WX6560,WX6561);
	or 	XG15911 	(WX6577,WX6574,WX6575);
	or 	XG15912 	(WX6591,WX6588,WX6589);
	or 	XG15913 	(WX6605,WX6602,WX6603);
	or 	XG15914 	(WX6619,WX6616,WX6617);
	or 	XG15915 	(WX6633,WX6630,WX6631);
	or 	XG15916 	(WX6647,WX6644,WX6645);
	or 	XG15917 	(WX6661,WX6658,WX6659);
	or 	XG15918 	(WX6675,WX6672,WX6673);
	or 	XG15919 	(WX6689,WX6686,WX6687);
	or 	XG15920 	(WX6703,WX6700,WX6701);
	or 	XG15921 	(WX6717,WX6714,WX6715);
	or 	XG15922 	(WX6731,WX6728,WX6729);
	or 	XG15923 	(WX6745,WX6742,WX6743);
	or 	XG15924 	(WX6759,WX6756,WX6757);
	or 	XG15925 	(WX6773,WX6770,WX6771);
	or 	XG15926 	(WX6787,WX6784,WX6785);
	or 	XG15927 	(WX6801,WX6798,WX6799);
	or 	XG15928 	(WX6815,WX6812,WX6813);
	or 	XG15929 	(WX6829,WX6826,WX6827);
	or 	XG15930 	(WX6843,WX6840,WX6841);
	or 	XG15931 	(WX6857,WX6854,WX6855);
	or 	XG15932 	(WX6871,WX6868,WX6869);
	or 	XG15933 	(WX6885,WX6882,WX6883);
	or 	XG15934 	(WX6899,WX6896,WX6897);
	or 	XG15935 	(WX6913,WX6910,WX6911);
	or 	XG15936 	(WX6927,WX6924,WX6925);
	or 	XG15937 	(WX6941,WX6938,WX6939);
	or 	XG15938 	(WX5214,WX5211,WX5212);
	or 	XG15939 	(WX5228,WX5225,WX5226);
	or 	XG15940 	(WX5242,WX5239,WX5240);
	or 	XG15941 	(WX5256,WX5253,WX5254);
	or 	XG15942 	(WX5270,WX5267,WX5268);
	or 	XG15943 	(WX5284,WX5281,WX5282);
	or 	XG15944 	(WX5298,WX5295,WX5296);
	or 	XG15945 	(WX5312,WX5309,WX5310);
	or 	XG15946 	(WX5326,WX5323,WX5324);
	or 	XG15947 	(WX5340,WX5337,WX5338);
	or 	XG15948 	(WX5354,WX5351,WX5352);
	or 	XG15949 	(WX5368,WX5365,WX5366);
	or 	XG15950 	(WX5382,WX5379,WX5380);
	or 	XG15951 	(WX5396,WX5393,WX5394);
	or 	XG15952 	(WX5410,WX5407,WX5408);
	or 	XG15953 	(WX5424,WX5421,WX5422);
	or 	XG15954 	(WX5438,WX5435,WX5436);
	or 	XG15955 	(WX5452,WX5449,WX5450);
	or 	XG15956 	(WX5466,WX5463,WX5464);
	or 	XG15957 	(WX5480,WX5477,WX5478);
	or 	XG15958 	(WX5494,WX5491,WX5492);
	or 	XG15959 	(WX5508,WX5505,WX5506);
	or 	XG15960 	(WX5522,WX5519,WX5520);
	or 	XG15961 	(WX5536,WX5533,WX5534);
	or 	XG15962 	(WX5550,WX5547,WX5548);
	or 	XG15963 	(WX5564,WX5561,WX5562);
	or 	XG15964 	(WX5578,WX5575,WX5576);
	or 	XG15965 	(WX5592,WX5589,WX5590);
	or 	XG15966 	(WX5606,WX5603,WX5604);
	or 	XG15967 	(WX5620,WX5617,WX5618);
	or 	XG15968 	(WX5634,WX5631,WX5632);
	or 	XG15969 	(WX5648,WX5645,WX5646);
	or 	XG15970 	(WX3921,WX3918,WX3919);
	or 	XG15971 	(WX3935,WX3932,WX3933);
	or 	XG15972 	(WX3949,WX3946,WX3947);
	or 	XG15973 	(WX3963,WX3960,WX3961);
	or 	XG15974 	(WX3977,WX3974,WX3975);
	or 	XG15975 	(WX3991,WX3988,WX3989);
	or 	XG15976 	(WX4005,WX4002,WX4003);
	or 	XG15977 	(WX4019,WX4016,WX4017);
	or 	XG15978 	(WX4033,WX4030,WX4031);
	or 	XG15979 	(WX4047,WX4044,WX4045);
	or 	XG15980 	(WX4061,WX4058,WX4059);
	or 	XG15981 	(WX4075,WX4072,WX4073);
	or 	XG15982 	(WX4089,WX4086,WX4087);
	or 	XG15983 	(WX4103,WX4100,WX4101);
	or 	XG15984 	(WX4117,WX4114,WX4115);
	or 	XG15985 	(WX4131,WX4128,WX4129);
	or 	XG15986 	(WX4145,WX4142,WX4143);
	or 	XG15987 	(WX4159,WX4156,WX4157);
	or 	XG15988 	(WX4173,WX4170,WX4171);
	or 	XG15989 	(WX4187,WX4184,WX4185);
	or 	XG15990 	(WX4201,WX4198,WX4199);
	or 	XG15991 	(WX4215,WX4212,WX4213);
	or 	XG15992 	(WX4229,WX4226,WX4227);
	or 	XG15993 	(WX4243,WX4240,WX4241);
	or 	XG15994 	(WX4257,WX4254,WX4255);
	or 	XG15995 	(WX4271,WX4268,WX4269);
	or 	XG15996 	(WX4285,WX4282,WX4283);
	or 	XG15997 	(WX4299,WX4296,WX4297);
	or 	XG15998 	(WX4313,WX4310,WX4311);
	or 	XG15999 	(WX4327,WX4324,WX4325);
	or 	XG16000 	(WX4341,WX4338,WX4339);
	or 	XG16001 	(WX4355,WX4352,WX4353);
	or 	XG16002 	(WX2628,WX2625,WX2626);
	or 	XG16003 	(WX2642,WX2639,WX2640);
	or 	XG16004 	(WX2656,WX2653,WX2654);
	or 	XG16005 	(WX2670,WX2667,WX2668);
	or 	XG16006 	(WX2684,WX2681,WX2682);
	or 	XG16007 	(WX2698,WX2695,WX2696);
	or 	XG16008 	(WX2712,WX2709,WX2710);
	or 	XG16009 	(WX2726,WX2723,WX2724);
	or 	XG16010 	(WX2740,WX2737,WX2738);
	or 	XG16011 	(WX2754,WX2751,WX2752);
	or 	XG16012 	(WX2768,WX2765,WX2766);
	or 	XG16013 	(WX2782,WX2779,WX2780);
	or 	XG16014 	(WX2796,WX2793,WX2794);
	or 	XG16015 	(WX2810,WX2807,WX2808);
	or 	XG16016 	(WX2824,WX2821,WX2822);
	or 	XG16017 	(WX2838,WX2835,WX2836);
	or 	XG16018 	(WX2852,WX2849,WX2850);
	or 	XG16019 	(WX2866,WX2863,WX2864);
	or 	XG16020 	(WX2880,WX2877,WX2878);
	or 	XG16021 	(WX2894,WX2891,WX2892);
	or 	XG16022 	(WX2908,WX2905,WX2906);
	or 	XG16023 	(WX2922,WX2919,WX2920);
	or 	XG16024 	(WX2936,WX2933,WX2934);
	or 	XG16025 	(WX2950,WX2947,WX2948);
	or 	XG16026 	(WX2964,WX2961,WX2962);
	or 	XG16027 	(WX2978,WX2975,WX2976);
	or 	XG16028 	(WX2992,WX2989,WX2990);
	or 	XG16029 	(WX3006,WX3003,WX3004);
	or 	XG16030 	(WX3020,WX3017,WX3018);
	or 	XG16031 	(WX3034,WX3031,WX3032);
	or 	XG16032 	(WX3048,WX3045,WX3046);
	or 	XG16033 	(WX3062,WX3059,WX3060);
	or 	XG16034 	(WX1335,WX1332,WX1333);
	or 	XG16035 	(WX1349,WX1346,WX1347);
	or 	XG16036 	(WX1363,WX1360,WX1361);
	or 	XG16037 	(WX1377,WX1374,WX1375);
	or 	XG16038 	(WX1391,WX1388,WX1389);
	or 	XG16039 	(WX1405,WX1402,WX1403);
	or 	XG16040 	(WX1419,WX1416,WX1417);
	or 	XG16041 	(WX1433,WX1430,WX1431);
	or 	XG16042 	(WX1447,WX1444,WX1445);
	or 	XG16043 	(WX1461,WX1458,WX1459);
	or 	XG16044 	(WX1475,WX1472,WX1473);
	or 	XG16045 	(WX1489,WX1486,WX1487);
	or 	XG16046 	(WX1503,WX1500,WX1501);
	or 	XG16047 	(WX1517,WX1514,WX1515);
	or 	XG16048 	(WX1531,WX1528,WX1529);
	or 	XG16049 	(WX1545,WX1542,WX1543);
	or 	XG16050 	(WX1559,WX1556,WX1557);
	or 	XG16051 	(WX1573,WX1570,WX1571);
	or 	XG16052 	(WX1587,WX1584,WX1585);
	or 	XG16053 	(WX1601,WX1598,WX1599);
	or 	XG16054 	(WX1615,WX1612,WX1613);
	or 	XG16055 	(WX1629,WX1626,WX1627);
	or 	XG16056 	(WX1643,WX1640,WX1641);
	or 	XG16057 	(WX1657,WX1654,WX1655);
	or 	XG16058 	(WX1671,WX1668,WX1669);
	or 	XG16059 	(WX1685,WX1682,WX1683);
	or 	XG16060 	(WX1699,WX1696,WX1697);
	or 	XG16061 	(WX1713,WX1710,WX1711);
	or 	XG16062 	(WX1727,WX1724,WX1725);
	or 	XG16063 	(WX1741,WX1738,WX1739);
	or 	XG16064 	(WX1755,WX1752,WX1753);
	or 	XG16065 	(WX1769,WX1766,WX1767);
	or 	XG16066 	(WX42,WX39,WX40);
	or 	XG16067 	(WX56,WX53,WX54);
	or 	XG16068 	(WX70,WX67,WX68);
	or 	XG16069 	(WX84,WX81,WX82);
	or 	XG16070 	(WX98,WX95,WX96);
	or 	XG16071 	(WX112,WX109,WX110);
	or 	XG16072 	(WX126,WX123,WX124);
	or 	XG16073 	(WX140,WX137,WX138);
	or 	XG16074 	(WX154,WX151,WX152);
	or 	XG16075 	(WX168,WX165,WX166);
	or 	XG16076 	(WX182,WX179,WX180);
	or 	XG16077 	(WX196,WX193,WX194);
	or 	XG16078 	(WX210,WX207,WX208);
	or 	XG16079 	(WX224,WX221,WX222);
	or 	XG16080 	(WX238,WX235,WX236);
	or 	XG16081 	(WX252,WX249,WX250);
	or 	XG16082 	(WX266,WX263,WX264);
	or 	XG16083 	(WX280,WX277,WX278);
	or 	XG16084 	(WX294,WX291,WX292);
	or 	XG16085 	(WX308,WX305,WX306);
	or 	XG16086 	(WX322,WX319,WX320);
	or 	XG16087 	(WX336,WX333,WX334);
	or 	XG16088 	(WX350,WX347,WX348);
	or 	XG16089 	(WX364,WX361,WX362);
	or 	XG16090 	(WX378,WX375,WX376);
	or 	XG16091 	(WX392,WX389,WX390);
	or 	XG16092 	(WX406,WX403,WX404);
	or 	XG16093 	(WX420,WX417,WX418);
	or 	XG16094 	(WX434,WX431,WX432);
	or 	XG16095 	(WX448,WX445,WX446);
	or 	XG16096 	(WX462,WX459,WX460);
	or 	XG16097 	(WX476,WX473,WX474);
	and 	XG16098 	(WX10813,WX11347,WX10824);
	and 	XG16099 	(WX10799,WX11347,WX10810);
	and 	XG16100 	(WX10785,WX11347,WX10796);
	and 	XG16101 	(WX10771,WX11347,WX10782);
	and 	XG16102 	(WX10757,WX11347,WX10768);
	and 	XG16103 	(WX10743,WX11347,WX10754);
	and 	XG16104 	(WX10729,WX11347,WX10740);
	and 	XG16105 	(WX10715,WX11347,WX10726);
	and 	XG16106 	(WX10701,WX11347,WX10712);
	and 	XG16107 	(WX10687,WX11347,WX10698);
	and 	XG16108 	(WX10673,WX11347,WX10684);
	and 	XG16109 	(WX10659,WX11347,WX10670);
	and 	XG16110 	(WX10645,WX11347,WX10656);
	and 	XG16111 	(WX10631,WX11347,WX10642);
	and 	XG16112 	(WX10617,WX11347,WX10628);
	and 	XG16113 	(WX10603,WX11347,WX10614);
	and 	XG16114 	(WX10589,WX11347,WX10600);
	and 	XG16115 	(WX10575,WX11347,WX10586);
	and 	XG16116 	(WX10561,WX11347,WX10572);
	and 	XG16117 	(WX10547,WX11347,WX10558);
	and 	XG16118 	(WX10533,WX11347,WX10544);
	and 	XG16119 	(WX10519,WX11347,WX10530);
	and 	XG16120 	(WX10505,WX11347,WX10516);
	and 	XG16121 	(WX10491,WX11347,WX10502);
	and 	XG16122 	(WX10477,WX11347,WX10488);
	and 	XG16123 	(WX10463,WX11347,WX10474);
	and 	XG16124 	(WX10449,WX11347,WX10460);
	and 	XG16125 	(WX10435,WX11347,WX10446);
	and 	XG16126 	(WX10421,WX11347,WX10432);
	and 	XG16127 	(WX10407,WX11347,WX10418);
	and 	XG16128 	(WX10393,WX11347,WX10404);
	and 	XG16129 	(WX10379,WX11347,WX10390);
	and 	XG16130 	(WX9520,WX10054,WX9531);
	and 	XG16131 	(WX9506,WX10054,WX9517);
	and 	XG16132 	(WX9492,WX10054,WX9503);
	and 	XG16133 	(WX9478,WX10054,WX9489);
	and 	XG16134 	(WX9464,WX10054,WX9475);
	and 	XG16135 	(WX9450,WX10054,WX9461);
	and 	XG16136 	(WX9436,WX10054,WX9447);
	and 	XG16137 	(WX9422,WX10054,WX9433);
	and 	XG16138 	(WX9408,WX10054,WX9419);
	and 	XG16139 	(WX9394,WX10054,WX9405);
	and 	XG16140 	(WX9380,WX10054,WX9391);
	and 	XG16141 	(WX9366,WX10054,WX9377);
	and 	XG16142 	(WX9352,WX10054,WX9363);
	and 	XG16143 	(WX9338,WX10054,WX9349);
	and 	XG16144 	(WX9324,WX10054,WX9335);
	and 	XG16145 	(WX9310,WX10054,WX9321);
	and 	XG16146 	(WX9296,WX10054,WX9307);
	and 	XG16147 	(WX9282,WX10054,WX9293);
	and 	XG16148 	(WX9268,WX10054,WX9279);
	and 	XG16149 	(WX9254,WX10054,WX9265);
	and 	XG16150 	(WX9240,WX10054,WX9251);
	and 	XG16151 	(WX9226,WX10054,WX9237);
	and 	XG16152 	(WX9212,WX10054,WX9223);
	and 	XG16153 	(WX9198,WX10054,WX9209);
	and 	XG16154 	(WX9184,WX10054,WX9195);
	and 	XG16155 	(WX9170,WX10054,WX9181);
	and 	XG16156 	(WX9156,WX10054,WX9167);
	and 	XG16157 	(WX9142,WX10054,WX9153);
	and 	XG16158 	(WX9128,WX10054,WX9139);
	and 	XG16159 	(WX9114,WX10054,WX9125);
	and 	XG16160 	(WX9100,WX10054,WX9111);
	and 	XG16161 	(WX9086,WX10054,WX9097);
	and 	XG16162 	(WX8227,WX8761,WX8238);
	and 	XG16163 	(WX8213,WX8761,WX8224);
	and 	XG16164 	(WX8199,WX8761,WX8210);
	and 	XG16165 	(WX8185,WX8761,WX8196);
	and 	XG16166 	(WX8171,WX8761,WX8182);
	and 	XG16167 	(WX8157,WX8761,WX8168);
	and 	XG16168 	(WX8143,WX8761,WX8154);
	and 	XG16169 	(WX8129,WX8761,WX8140);
	and 	XG16170 	(WX8115,WX8761,WX8126);
	and 	XG16171 	(WX8101,WX8761,WX8112);
	and 	XG16172 	(WX8087,WX8761,WX8098);
	and 	XG16173 	(WX8073,WX8761,WX8084);
	and 	XG16174 	(WX8059,WX8761,WX8070);
	and 	XG16175 	(WX8045,WX8761,WX8056);
	and 	XG16176 	(WX8031,WX8761,WX8042);
	and 	XG16177 	(WX8017,WX8761,WX8028);
	and 	XG16178 	(WX8003,WX8761,WX8014);
	and 	XG16179 	(WX7989,WX8761,WX8000);
	and 	XG16180 	(WX7975,WX8761,WX7986);
	and 	XG16181 	(WX7961,WX8761,WX7972);
	and 	XG16182 	(WX7947,WX8761,WX7958);
	and 	XG16183 	(WX7933,WX8761,WX7944);
	and 	XG16184 	(WX7919,WX8761,WX7930);
	and 	XG16185 	(WX7905,WX8761,WX7916);
	and 	XG16186 	(WX7891,WX8761,WX7902);
	and 	XG16187 	(WX7877,WX8761,WX7888);
	and 	XG16188 	(WX7863,WX8761,WX7874);
	and 	XG16189 	(WX7849,WX8761,WX7860);
	and 	XG16190 	(WX7835,WX8761,WX7846);
	and 	XG16191 	(WX7821,WX8761,WX7832);
	and 	XG16192 	(WX7807,WX8761,WX7818);
	and 	XG16193 	(WX7793,WX8761,WX7804);
	and 	XG16194 	(WX6934,WX7468,WX6945);
	and 	XG16195 	(WX6920,WX7468,WX6931);
	and 	XG16196 	(WX6906,WX7468,WX6917);
	and 	XG16197 	(WX6892,WX7468,WX6903);
	and 	XG16198 	(WX6878,WX7468,WX6889);
	and 	XG16199 	(WX6864,WX7468,WX6875);
	and 	XG16200 	(WX6850,WX7468,WX6861);
	and 	XG16201 	(WX6836,WX7468,WX6847);
	and 	XG16202 	(WX6822,WX7468,WX6833);
	and 	XG16203 	(WX6808,WX7468,WX6819);
	and 	XG16204 	(WX6794,WX7468,WX6805);
	and 	XG16205 	(WX6780,WX7468,WX6791);
	and 	XG16206 	(WX6766,WX7468,WX6777);
	and 	XG16207 	(WX6752,WX7468,WX6763);
	and 	XG16208 	(WX6738,WX7468,WX6749);
	and 	XG16209 	(WX6724,WX7468,WX6735);
	and 	XG16210 	(WX6710,WX7468,WX6721);
	and 	XG16211 	(WX6696,WX7468,WX6707);
	and 	XG16212 	(WX6682,WX7468,WX6693);
	and 	XG16213 	(WX6668,WX7468,WX6679);
	and 	XG16214 	(WX6654,WX7468,WX6665);
	and 	XG16215 	(WX6640,WX7468,WX6651);
	and 	XG16216 	(WX6626,WX7468,WX6637);
	and 	XG16217 	(WX6612,WX7468,WX6623);
	and 	XG16218 	(WX6598,WX7468,WX6609);
	and 	XG16219 	(WX6584,WX7468,WX6595);
	and 	XG16220 	(WX6570,WX7468,WX6581);
	and 	XG16221 	(WX6556,WX7468,WX6567);
	and 	XG16222 	(WX6542,WX7468,WX6553);
	and 	XG16223 	(WX6528,WX7468,WX6539);
	and 	XG16224 	(WX6514,WX7468,WX6525);
	and 	XG16225 	(WX6500,WX7468,WX6511);
	and 	XG16226 	(WX5641,WX6175,WX5652);
	and 	XG16227 	(WX5627,WX6175,WX5638);
	and 	XG16228 	(WX5613,WX6175,WX5624);
	and 	XG16229 	(WX5599,WX6175,WX5610);
	and 	XG16230 	(WX5585,WX6175,WX5596);
	and 	XG16231 	(WX5571,WX6175,WX5582);
	and 	XG16232 	(WX5557,WX6175,WX5568);
	and 	XG16233 	(WX5543,WX6175,WX5554);
	and 	XG16234 	(WX5529,WX6175,WX5540);
	and 	XG16235 	(WX5515,WX6175,WX5526);
	and 	XG16236 	(WX5501,WX6175,WX5512);
	and 	XG16237 	(WX5487,WX6175,WX5498);
	and 	XG16238 	(WX5473,WX6175,WX5484);
	and 	XG16239 	(WX5459,WX6175,WX5470);
	and 	XG16240 	(WX5445,WX6175,WX5456);
	and 	XG16241 	(WX5431,WX6175,WX5442);
	and 	XG16242 	(WX5417,WX6175,WX5428);
	and 	XG16243 	(WX5403,WX6175,WX5414);
	and 	XG16244 	(WX5389,WX6175,WX5400);
	and 	XG16245 	(WX5375,WX6175,WX5386);
	and 	XG16246 	(WX5361,WX6175,WX5372);
	and 	XG16247 	(WX5347,WX6175,WX5358);
	and 	XG16248 	(WX5333,WX6175,WX5344);
	and 	XG16249 	(WX5319,WX6175,WX5330);
	and 	XG16250 	(WX5305,WX6175,WX5316);
	and 	XG16251 	(WX5291,WX6175,WX5302);
	and 	XG16252 	(WX5277,WX6175,WX5288);
	and 	XG16253 	(WX5263,WX6175,WX5274);
	and 	XG16254 	(WX5249,WX6175,WX5260);
	and 	XG16255 	(WX5235,WX6175,WX5246);
	and 	XG16256 	(WX5221,WX6175,WX5232);
	and 	XG16257 	(WX5207,WX6175,WX5218);
	and 	XG16258 	(WX4348,WX4882,WX4359);
	and 	XG16259 	(WX4334,WX4882,WX4345);
	and 	XG16260 	(WX4320,WX4882,WX4331);
	and 	XG16261 	(WX4306,WX4882,WX4317);
	and 	XG16262 	(WX4292,WX4882,WX4303);
	and 	XG16263 	(WX4278,WX4882,WX4289);
	and 	XG16264 	(WX4264,WX4882,WX4275);
	and 	XG16265 	(WX4250,WX4882,WX4261);
	and 	XG16266 	(WX4236,WX4882,WX4247);
	and 	XG16267 	(WX4222,WX4882,WX4233);
	and 	XG16268 	(WX4208,WX4882,WX4219);
	and 	XG16269 	(WX4194,WX4882,WX4205);
	and 	XG16270 	(WX4180,WX4882,WX4191);
	and 	XG16271 	(WX4166,WX4882,WX4177);
	and 	XG16272 	(WX4152,WX4882,WX4163);
	and 	XG16273 	(WX4138,WX4882,WX4149);
	and 	XG16274 	(WX4124,WX4882,WX4135);
	and 	XG16275 	(WX4110,WX4882,WX4121);
	and 	XG16276 	(WX4096,WX4882,WX4107);
	and 	XG16277 	(WX4082,WX4882,WX4093);
	and 	XG16278 	(WX4068,WX4882,WX4079);
	and 	XG16279 	(WX4054,WX4882,WX4065);
	and 	XG16280 	(WX4040,WX4882,WX4051);
	and 	XG16281 	(WX4026,WX4882,WX4037);
	and 	XG16282 	(WX4012,WX4882,WX4023);
	and 	XG16283 	(WX3998,WX4882,WX4009);
	and 	XG16284 	(WX3984,WX4882,WX3995);
	and 	XG16285 	(WX3970,WX4882,WX3981);
	and 	XG16286 	(WX3956,WX4882,WX3967);
	and 	XG16287 	(WX3942,WX4882,WX3953);
	and 	XG16288 	(WX3928,WX4882,WX3939);
	and 	XG16289 	(WX3914,WX4882,WX3925);
	and 	XG16290 	(WX3055,WX3589,WX3066);
	and 	XG16291 	(WX3041,WX3589,WX3052);
	and 	XG16292 	(WX3027,WX3589,WX3038);
	and 	XG16293 	(WX3013,WX3589,WX3024);
	and 	XG16294 	(WX2999,WX3589,WX3010);
	and 	XG16295 	(WX2985,WX3589,WX2996);
	and 	XG16296 	(WX2971,WX3589,WX2982);
	and 	XG16297 	(WX2957,WX3589,WX2968);
	and 	XG16298 	(WX2943,WX3589,WX2954);
	and 	XG16299 	(WX2929,WX3589,WX2940);
	and 	XG16300 	(WX2915,WX3589,WX2926);
	and 	XG16301 	(WX2901,WX3589,WX2912);
	and 	XG16302 	(WX2887,WX3589,WX2898);
	and 	XG16303 	(WX2873,WX3589,WX2884);
	and 	XG16304 	(WX2859,WX3589,WX2870);
	and 	XG16305 	(WX2845,WX3589,WX2856);
	and 	XG16306 	(WX2831,WX3589,WX2842);
	and 	XG16307 	(WX2817,WX3589,WX2828);
	and 	XG16308 	(WX2803,WX3589,WX2814);
	and 	XG16309 	(WX2789,WX3589,WX2800);
	and 	XG16310 	(WX2775,WX3589,WX2786);
	and 	XG16311 	(WX2761,WX3589,WX2772);
	and 	XG16312 	(WX2747,WX3589,WX2758);
	and 	XG16313 	(WX2733,WX3589,WX2744);
	and 	XG16314 	(WX2719,WX3589,WX2730);
	and 	XG16315 	(WX2705,WX3589,WX2716);
	and 	XG16316 	(WX2691,WX3589,WX2702);
	and 	XG16317 	(WX2677,WX3589,WX2688);
	and 	XG16318 	(WX2663,WX3589,WX2674);
	and 	XG16319 	(WX2649,WX3589,WX2660);
	and 	XG16320 	(WX2635,WX3589,WX2646);
	and 	XG16321 	(WX2621,WX3589,WX2632);
	and 	XG16322 	(WX1762,WX2296,WX1773);
	and 	XG16323 	(WX1748,WX2296,WX1759);
	and 	XG16324 	(WX1734,WX2296,WX1745);
	and 	XG16325 	(WX1720,WX2296,WX1731);
	and 	XG16326 	(WX1706,WX2296,WX1717);
	and 	XG16327 	(WX1692,WX2296,WX1703);
	and 	XG16328 	(WX1678,WX2296,WX1689);
	and 	XG16329 	(WX1664,WX2296,WX1675);
	and 	XG16330 	(WX1650,WX2296,WX1661);
	and 	XG16331 	(WX1636,WX2296,WX1647);
	and 	XG16332 	(WX1622,WX2296,WX1633);
	and 	XG16333 	(WX1608,WX2296,WX1619);
	and 	XG16334 	(WX1594,WX2296,WX1605);
	and 	XG16335 	(WX1580,WX2296,WX1591);
	and 	XG16336 	(WX1566,WX2296,WX1577);
	and 	XG16337 	(WX1552,WX2296,WX1563);
	and 	XG16338 	(WX1538,WX2296,WX1549);
	and 	XG16339 	(WX1524,WX2296,WX1535);
	and 	XG16340 	(WX1510,WX2296,WX1521);
	and 	XG16341 	(WX1496,WX2296,WX1507);
	and 	XG16342 	(WX1482,WX2296,WX1493);
	and 	XG16343 	(WX1468,WX2296,WX1479);
	and 	XG16344 	(WX1454,WX2296,WX1465);
	and 	XG16345 	(WX1440,WX2296,WX1451);
	and 	XG16346 	(WX1426,WX2296,WX1437);
	and 	XG16347 	(WX1412,WX2296,WX1423);
	and 	XG16348 	(WX1398,WX2296,WX1409);
	and 	XG16349 	(WX1384,WX2296,WX1395);
	and 	XG16350 	(WX1370,WX2296,WX1381);
	and 	XG16351 	(WX1356,WX2296,WX1367);
	and 	XG16352 	(WX1342,WX2296,WX1353);
	and 	XG16353 	(WX1328,WX2296,WX1339);
	and 	XG16354 	(WX469,WX1003,WX480);
	and 	XG16355 	(WX455,WX1003,WX466);
	and 	XG16356 	(WX441,WX1003,WX452);
	and 	XG16357 	(WX427,WX1003,WX438);
	and 	XG16358 	(WX413,WX1003,WX424);
	and 	XG16359 	(WX399,WX1003,WX410);
	and 	XG16360 	(WX385,WX1003,WX396);
	and 	XG16361 	(WX371,WX1003,WX382);
	and 	XG16362 	(WX357,WX1003,WX368);
	and 	XG16363 	(WX343,WX1003,WX354);
	and 	XG16364 	(WX329,WX1003,WX340);
	and 	XG16365 	(WX315,WX1003,WX326);
	and 	XG16366 	(WX301,WX1003,WX312);
	and 	XG16367 	(WX287,WX1003,WX298);
	and 	XG16368 	(WX273,WX1003,WX284);
	and 	XG16369 	(WX259,WX1003,WX270);
	and 	XG16370 	(WX245,WX1003,WX256);
	and 	XG16371 	(WX231,WX1003,WX242);
	and 	XG16372 	(WX217,WX1003,WX228);
	and 	XG16373 	(WX203,WX1003,WX214);
	and 	XG16374 	(WX189,WX1003,WX200);
	and 	XG16375 	(WX175,WX1003,WX186);
	and 	XG16376 	(WX161,WX1003,WX172);
	and 	XG16377 	(WX147,WX1003,WX158);
	and 	XG16378 	(WX133,WX1003,WX144);
	and 	XG16379 	(WX119,WX1003,WX130);
	and 	XG16380 	(WX105,WX1003,WX116);
	and 	XG16381 	(WX91,WX1003,WX102);
	and 	XG16382 	(WX77,WX1003,WX88);
	and 	XG16383 	(WX63,WX1003,WX74);
	and 	XG16384 	(WX49,WX1003,WX60);
	and 	XG16385 	(WX35,WX1003,WX46);
	and 	XG16386 	(WX9521,WX9522,WX9527);
	and 	XG16387 	(WX9507,WX9508,WX9513);
	and 	XG16388 	(WX9493,WX9494,WX9499);
	and 	XG16389 	(WX9479,WX9480,WX9485);
	and 	XG16390 	(WX9465,WX9466,WX9471);
	and 	XG16391 	(WX9451,WX9452,WX9457);
	and 	XG16392 	(WX9437,WX9438,WX9443);
	and 	XG16393 	(WX9423,WX9424,WX9429);
	and 	XG16394 	(WX9409,WX9410,WX9415);
	and 	XG16395 	(WX9395,WX9396,WX9401);
	and 	XG16396 	(WX9381,WX9382,WX9387);
	and 	XG16397 	(WX9367,WX9368,WX9373);
	and 	XG16398 	(WX9353,WX9354,WX9359);
	and 	XG16399 	(WX9339,WX9340,WX9345);
	and 	XG16400 	(WX9325,WX9326,WX9331);
	and 	XG16401 	(WX9311,WX9312,WX9317);
	and 	XG16402 	(WX9297,WX9298,WX9303);
	and 	XG16403 	(WX9283,WX9284,WX9289);
	and 	XG16404 	(WX9269,WX9270,WX9275);
	and 	XG16405 	(WX9255,WX9256,WX9261);
	and 	XG16406 	(WX9241,WX9242,WX9247);
	and 	XG16407 	(WX9227,WX9228,WX9233);
	and 	XG16408 	(WX9213,WX9214,WX9219);
	and 	XG16409 	(WX9199,WX9200,WX9205);
	and 	XG16410 	(WX9185,WX9186,WX9191);
	and 	XG16411 	(WX9171,WX9172,WX9177);
	and 	XG16412 	(WX9157,WX9158,WX9163);
	and 	XG16413 	(WX9143,WX9144,WX9149);
	and 	XG16414 	(WX9129,WX9130,WX9135);
	and 	XG16415 	(WX9115,WX9116,WX9121);
	and 	XG16416 	(WX9101,WX9102,WX9107);
	and 	XG16417 	(WX9087,WX9088,WX9093);
	and 	XG16418 	(WX8228,WX8229,WX8234);
	and 	XG16419 	(WX8214,WX8215,WX8220);
	and 	XG16420 	(WX8200,WX8201,WX8206);
	and 	XG16421 	(WX8186,WX8187,WX8192);
	and 	XG16422 	(WX8172,WX8173,WX8178);
	and 	XG16423 	(WX8158,WX8159,WX8164);
	and 	XG16424 	(WX8144,WX8145,WX8150);
	and 	XG16425 	(WX8130,WX8131,WX8136);
	and 	XG16426 	(WX8116,WX8117,WX8122);
	and 	XG16427 	(WX8102,WX8103,WX8108);
	and 	XG16428 	(WX8088,WX8089,WX8094);
	and 	XG16429 	(WX8074,WX8075,WX8080);
	and 	XG16430 	(WX8060,WX8061,WX8066);
	and 	XG16431 	(WX8046,WX8047,WX8052);
	and 	XG16432 	(WX8032,WX8033,WX8038);
	and 	XG16433 	(WX8018,WX8019,WX8024);
	and 	XG16434 	(WX8004,WX8005,WX8010);
	and 	XG16435 	(WX7990,WX7991,WX7996);
	and 	XG16436 	(WX7976,WX7977,WX7982);
	and 	XG16437 	(WX7962,WX7963,WX7968);
	and 	XG16438 	(WX7948,WX7949,WX7954);
	and 	XG16439 	(WX7934,WX7935,WX7940);
	and 	XG16440 	(WX7920,WX7921,WX7926);
	and 	XG16441 	(WX7906,WX7907,WX7912);
	and 	XG16442 	(WX7892,WX7893,WX7898);
	and 	XG16443 	(WX7878,WX7879,WX7884);
	and 	XG16444 	(WX7864,WX7865,WX7870);
	and 	XG16445 	(WX7850,WX7851,WX7856);
	and 	XG16446 	(WX7836,WX7837,WX7842);
	and 	XG16447 	(WX7822,WX7823,WX7828);
	and 	XG16448 	(WX7808,WX7809,WX7814);
	and 	XG16449 	(WX7794,WX7795,WX7800);
	and 	XG16450 	(WX6935,WX6936,WX6941);
	and 	XG16451 	(WX6921,WX6922,WX6927);
	and 	XG16452 	(WX6907,WX6908,WX6913);
	and 	XG16453 	(WX6893,WX6894,WX6899);
	and 	XG16454 	(WX6879,WX6880,WX6885);
	and 	XG16455 	(WX6865,WX6866,WX6871);
	and 	XG16456 	(WX6851,WX6852,WX6857);
	and 	XG16457 	(WX6837,WX6838,WX6843);
	and 	XG16458 	(WX6823,WX6824,WX6829);
	and 	XG16459 	(WX6809,WX6810,WX6815);
	and 	XG16460 	(WX6795,WX6796,WX6801);
	and 	XG16461 	(WX6781,WX6782,WX6787);
	and 	XG16462 	(WX6767,WX6768,WX6773);
	and 	XG16463 	(WX6753,WX6754,WX6759);
	and 	XG16464 	(WX6739,WX6740,WX6745);
	and 	XG16465 	(WX6725,WX6726,WX6731);
	and 	XG16466 	(WX6711,WX6712,WX6717);
	and 	XG16467 	(WX6697,WX6698,WX6703);
	and 	XG16468 	(WX6683,WX6684,WX6689);
	and 	XG16469 	(WX6669,WX6670,WX6675);
	and 	XG16470 	(WX6655,WX6656,WX6661);
	and 	XG16471 	(WX6641,WX6642,WX6647);
	and 	XG16472 	(WX6627,WX6628,WX6633);
	and 	XG16473 	(WX6613,WX6614,WX6619);
	and 	XG16474 	(WX6599,WX6600,WX6605);
	and 	XG16475 	(WX6585,WX6586,WX6591);
	and 	XG16476 	(WX6571,WX6572,WX6577);
	and 	XG16477 	(WX6557,WX6558,WX6563);
	and 	XG16478 	(WX6543,WX6544,WX6549);
	and 	XG16479 	(WX6529,WX6530,WX6535);
	and 	XG16480 	(WX6515,WX6516,WX6521);
	and 	XG16481 	(WX6501,WX6502,WX6507);
	and 	XG16482 	(WX5642,WX5643,WX5648);
	and 	XG16483 	(WX5628,WX5629,WX5634);
	and 	XG16484 	(WX5614,WX5615,WX5620);
	and 	XG16485 	(WX5600,WX5601,WX5606);
	and 	XG16486 	(WX5586,WX5587,WX5592);
	and 	XG16487 	(WX5572,WX5573,WX5578);
	and 	XG16488 	(WX5558,WX5559,WX5564);
	and 	XG16489 	(WX5544,WX5545,WX5550);
	and 	XG16490 	(WX5530,WX5531,WX5536);
	and 	XG16491 	(WX5516,WX5517,WX5522);
	and 	XG16492 	(WX5502,WX5503,WX5508);
	and 	XG16493 	(WX5488,WX5489,WX5494);
	and 	XG16494 	(WX5474,WX5475,WX5480);
	and 	XG16495 	(WX5460,WX5461,WX5466);
	and 	XG16496 	(WX5446,WX5447,WX5452);
	and 	XG16497 	(WX5432,WX5433,WX5438);
	and 	XG16498 	(WX5418,WX5419,WX5424);
	and 	XG16499 	(WX5404,WX5405,WX5410);
	and 	XG16500 	(WX5390,WX5391,WX5396);
	and 	XG16501 	(WX5376,WX5377,WX5382);
	and 	XG16502 	(WX5362,WX5363,WX5368);
	and 	XG16503 	(WX5348,WX5349,WX5354);
	and 	XG16504 	(WX5334,WX5335,WX5340);
	and 	XG16505 	(WX5320,WX5321,WX5326);
	and 	XG16506 	(WX5306,WX5307,WX5312);
	and 	XG16507 	(WX5292,WX5293,WX5298);
	and 	XG16508 	(WX5278,WX5279,WX5284);
	and 	XG16509 	(WX5264,WX5265,WX5270);
	and 	XG16510 	(WX5250,WX5251,WX5256);
	and 	XG16511 	(WX5236,WX5237,WX5242);
	and 	XG16512 	(WX5222,WX5223,WX5228);
	and 	XG16513 	(WX5208,WX5209,WX5214);
	and 	XG16514 	(WX4349,WX4350,WX4355);
	and 	XG16515 	(WX4335,WX4336,WX4341);
	and 	XG16516 	(WX4321,WX4322,WX4327);
	and 	XG16517 	(WX4307,WX4308,WX4313);
	and 	XG16518 	(WX4293,WX4294,WX4299);
	and 	XG16519 	(WX4279,WX4280,WX4285);
	and 	XG16520 	(WX4265,WX4266,WX4271);
	and 	XG16521 	(WX4251,WX4252,WX4257);
	and 	XG16522 	(WX4237,WX4238,WX4243);
	and 	XG16523 	(WX4223,WX4224,WX4229);
	and 	XG16524 	(WX4209,WX4210,WX4215);
	and 	XG16525 	(WX4195,WX4196,WX4201);
	and 	XG16526 	(WX4181,WX4182,WX4187);
	and 	XG16527 	(WX4167,WX4168,WX4173);
	and 	XG16528 	(WX4153,WX4154,WX4159);
	and 	XG16529 	(WX4139,WX4140,WX4145);
	and 	XG16530 	(WX4125,WX4126,WX4131);
	and 	XG16531 	(WX4111,WX4112,WX4117);
	and 	XG16532 	(WX4097,WX4098,WX4103);
	and 	XG16533 	(WX4083,WX4084,WX4089);
	and 	XG16534 	(WX4069,WX4070,WX4075);
	and 	XG16535 	(WX4055,WX4056,WX4061);
	and 	XG16536 	(WX4041,WX4042,WX4047);
	and 	XG16537 	(WX4027,WX4028,WX4033);
	and 	XG16538 	(WX4013,WX4014,WX4019);
	and 	XG16539 	(WX3999,WX4000,WX4005);
	and 	XG16540 	(WX3985,WX3986,WX3991);
	and 	XG16541 	(WX3971,WX3972,WX3977);
	and 	XG16542 	(WX3957,WX3958,WX3963);
	and 	XG16543 	(WX3943,WX3944,WX3949);
	and 	XG16544 	(WX3929,WX3930,WX3935);
	and 	XG16545 	(WX3915,WX3916,WX3921);
	and 	XG16546 	(WX3056,WX3057,WX3062);
	and 	XG16547 	(WX3042,WX3043,WX3048);
	and 	XG16548 	(WX3028,WX3029,WX3034);
	and 	XG16549 	(WX3014,WX3015,WX3020);
	and 	XG16550 	(WX3000,WX3001,WX3006);
	and 	XG16551 	(WX2986,WX2987,WX2992);
	and 	XG16552 	(WX2972,WX2973,WX2978);
	and 	XG16553 	(WX2958,WX2959,WX2964);
	and 	XG16554 	(WX2944,WX2945,WX2950);
	and 	XG16555 	(WX2930,WX2931,WX2936);
	and 	XG16556 	(WX2916,WX2917,WX2922);
	and 	XG16557 	(WX2902,WX2903,WX2908);
	and 	XG16558 	(WX2888,WX2889,WX2894);
	and 	XG16559 	(WX2874,WX2875,WX2880);
	and 	XG16560 	(WX2860,WX2861,WX2866);
	and 	XG16561 	(WX2846,WX2847,WX2852);
	and 	XG16562 	(WX2832,WX2833,WX2838);
	and 	XG16563 	(WX2818,WX2819,WX2824);
	and 	XG16564 	(WX2804,WX2805,WX2810);
	and 	XG16565 	(WX2790,WX2791,WX2796);
	and 	XG16566 	(WX2776,WX2777,WX2782);
	and 	XG16567 	(WX2762,WX2763,WX2768);
	and 	XG16568 	(WX2748,WX2749,WX2754);
	and 	XG16569 	(WX2734,WX2735,WX2740);
	and 	XG16570 	(WX2720,WX2721,WX2726);
	and 	XG16571 	(WX2706,WX2707,WX2712);
	and 	XG16572 	(WX2692,WX2693,WX2698);
	and 	XG16573 	(WX2678,WX2679,WX2684);
	and 	XG16574 	(WX2664,WX2665,WX2670);
	and 	XG16575 	(WX2650,WX2651,WX2656);
	and 	XG16576 	(WX2636,WX2637,WX2642);
	and 	XG16577 	(WX2622,WX2623,WX2628);
	and 	XG16578 	(WX1763,WX1764,WX1769);
	and 	XG16579 	(WX1749,WX1750,WX1755);
	and 	XG16580 	(WX1735,WX1736,WX1741);
	and 	XG16581 	(WX1721,WX1722,WX1727);
	and 	XG16582 	(WX1707,WX1708,WX1713);
	and 	XG16583 	(WX1693,WX1694,WX1699);
	and 	XG16584 	(WX1679,WX1680,WX1685);
	and 	XG16585 	(WX1665,WX1666,WX1671);
	and 	XG16586 	(WX1651,WX1652,WX1657);
	and 	XG16587 	(WX1637,WX1638,WX1643);
	and 	XG16588 	(WX1623,WX1624,WX1629);
	and 	XG16589 	(WX1609,WX1610,WX1615);
	and 	XG16590 	(WX1595,WX1596,WX1601);
	and 	XG16591 	(WX1581,WX1582,WX1587);
	and 	XG16592 	(WX1567,WX1568,WX1573);
	and 	XG16593 	(WX1553,WX1554,WX1559);
	and 	XG16594 	(WX1539,WX1540,WX1545);
	and 	XG16595 	(WX1525,WX1526,WX1531);
	and 	XG16596 	(WX1511,WX1512,WX1517);
	and 	XG16597 	(WX1497,WX1498,WX1503);
	and 	XG16598 	(WX1483,WX1484,WX1489);
	and 	XG16599 	(WX1469,WX1470,WX1475);
	and 	XG16600 	(WX1455,WX1456,WX1461);
	and 	XG16601 	(WX1441,WX1442,WX1447);
	and 	XG16602 	(WX1427,WX1428,WX1433);
	and 	XG16603 	(WX1413,WX1414,WX1419);
	and 	XG16604 	(WX1399,WX1400,WX1405);
	and 	XG16605 	(WX1385,WX1386,WX1391);
	and 	XG16606 	(WX1371,WX1372,WX1377);
	and 	XG16607 	(WX1357,WX1358,WX1363);
	and 	XG16608 	(WX1343,WX1344,WX1349);
	and 	XG16609 	(WX1329,WX1330,WX1335);
	and 	XG16610 	(WX470,WX471,WX476);
	and 	XG16611 	(WX456,WX457,WX462);
	and 	XG16612 	(WX442,WX443,WX448);
	and 	XG16613 	(WX428,WX429,WX434);
	and 	XG16614 	(WX414,WX415,WX420);
	and 	XG16615 	(WX400,WX401,WX406);
	and 	XG16616 	(WX386,WX387,WX392);
	and 	XG16617 	(WX372,WX373,WX378);
	and 	XG16618 	(WX358,WX359,WX364);
	and 	XG16619 	(WX344,WX345,WX350);
	and 	XG16620 	(WX330,WX331,WX336);
	and 	XG16621 	(WX316,WX317,WX322);
	and 	XG16622 	(WX302,WX303,WX308);
	and 	XG16623 	(WX288,WX289,WX294);
	and 	XG16624 	(WX274,WX275,WX280);
	and 	XG16625 	(WX260,WX261,WX266);
	and 	XG16626 	(WX246,WX247,WX252);
	and 	XG16627 	(WX232,WX233,WX238);
	and 	XG16628 	(WX218,WX219,WX224);
	and 	XG16629 	(WX204,WX205,WX210);
	and 	XG16630 	(WX190,WX191,WX196);
	and 	XG16631 	(WX176,WX177,WX182);
	and 	XG16632 	(WX162,WX163,WX168);
	and 	XG16633 	(WX148,WX149,WX154);
	and 	XG16634 	(WX134,WX135,WX140);
	and 	XG16635 	(WX120,WX121,WX126);
	and 	XG16636 	(WX106,WX107,WX112);
	and 	XG16637 	(WX92,WX93,WX98);
	and 	XG16638 	(WX78,WX79,WX84);
	and 	XG16639 	(WX64,WX65,WX70);
	and 	XG16640 	(WX50,WX51,WX56);
	and 	XG16641 	(WX36,WX37,WX42);
	or 	XG16642 	(WX38,WX35,WX36);
	or 	XG16643 	(WX52,WX49,WX50);
	or 	XG16644 	(WX66,WX63,WX64);
	or 	XG16645 	(WX80,WX77,WX78);
	or 	XG16646 	(WX94,WX91,WX92);
	or 	XG16647 	(WX108,WX105,WX106);
	or 	XG16648 	(WX122,WX119,WX120);
	or 	XG16649 	(WX136,WX133,WX134);
	or 	XG16650 	(WX150,WX147,WX148);
	or 	XG16651 	(WX164,WX161,WX162);
	or 	XG16652 	(WX178,WX175,WX176);
	or 	XG16653 	(WX192,WX189,WX190);
	or 	XG16654 	(WX206,WX203,WX204);
	or 	XG16655 	(WX220,WX217,WX218);
	or 	XG16656 	(WX234,WX231,WX232);
	or 	XG16657 	(WX248,WX245,WX246);
	or 	XG16658 	(WX262,WX259,WX260);
	or 	XG16659 	(WX276,WX273,WX274);
	or 	XG16660 	(WX290,WX287,WX288);
	or 	XG16661 	(WX304,WX301,WX302);
	or 	XG16662 	(WX318,WX315,WX316);
	or 	XG16663 	(WX332,WX329,WX330);
	or 	XG16664 	(WX346,WX343,WX344);
	or 	XG16665 	(WX360,WX357,WX358);
	or 	XG16666 	(WX374,WX371,WX372);
	or 	XG16667 	(WX388,WX385,WX386);
	or 	XG16668 	(WX402,WX399,WX400);
	or 	XG16669 	(WX416,WX413,WX414);
	or 	XG16670 	(WX430,WX427,WX428);
	or 	XG16671 	(WX444,WX441,WX442);
	or 	XG16672 	(WX458,WX455,WX456);
	or 	XG16673 	(WX472,WX469,WX470);
	or 	XG16674 	(WX1331,WX1328,WX1329);
	or 	XG16675 	(WX1345,WX1342,WX1343);
	or 	XG16676 	(WX1359,WX1356,WX1357);
	or 	XG16677 	(WX1373,WX1370,WX1371);
	or 	XG16678 	(WX1387,WX1384,WX1385);
	or 	XG16679 	(WX1401,WX1398,WX1399);
	or 	XG16680 	(WX1415,WX1412,WX1413);
	or 	XG16681 	(WX1429,WX1426,WX1427);
	or 	XG16682 	(WX1443,WX1440,WX1441);
	or 	XG16683 	(WX1457,WX1454,WX1455);
	or 	XG16684 	(WX1471,WX1468,WX1469);
	or 	XG16685 	(WX1485,WX1482,WX1483);
	or 	XG16686 	(WX1499,WX1496,WX1497);
	or 	XG16687 	(WX1513,WX1510,WX1511);
	or 	XG16688 	(WX1527,WX1524,WX1525);
	or 	XG16689 	(WX1541,WX1538,WX1539);
	or 	XG16690 	(WX1555,WX1552,WX1553);
	or 	XG16691 	(WX1569,WX1566,WX1567);
	or 	XG16692 	(WX1583,WX1580,WX1581);
	or 	XG16693 	(WX1597,WX1594,WX1595);
	or 	XG16694 	(WX1611,WX1608,WX1609);
	or 	XG16695 	(WX1625,WX1622,WX1623);
	or 	XG16696 	(WX1639,WX1636,WX1637);
	or 	XG16697 	(WX1653,WX1650,WX1651);
	or 	XG16698 	(WX1667,WX1664,WX1665);
	or 	XG16699 	(WX1681,WX1678,WX1679);
	or 	XG16700 	(WX1695,WX1692,WX1693);
	or 	XG16701 	(WX1709,WX1706,WX1707);
	or 	XG16702 	(WX1723,WX1720,WX1721);
	or 	XG16703 	(WX1737,WX1734,WX1735);
	or 	XG16704 	(WX1751,WX1748,WX1749);
	or 	XG16705 	(WX1765,WX1762,WX1763);
	or 	XG16706 	(WX2624,WX2621,WX2622);
	or 	XG16707 	(WX2638,WX2635,WX2636);
	or 	XG16708 	(WX2652,WX2649,WX2650);
	or 	XG16709 	(WX2666,WX2663,WX2664);
	or 	XG16710 	(WX2680,WX2677,WX2678);
	or 	XG16711 	(WX2694,WX2691,WX2692);
	or 	XG16712 	(WX2708,WX2705,WX2706);
	or 	XG16713 	(WX2722,WX2719,WX2720);
	or 	XG16714 	(WX2736,WX2733,WX2734);
	or 	XG16715 	(WX2750,WX2747,WX2748);
	or 	XG16716 	(WX2764,WX2761,WX2762);
	or 	XG16717 	(WX2778,WX2775,WX2776);
	or 	XG16718 	(WX2792,WX2789,WX2790);
	or 	XG16719 	(WX2806,WX2803,WX2804);
	or 	XG16720 	(WX2820,WX2817,WX2818);
	or 	XG16721 	(WX2834,WX2831,WX2832);
	or 	XG16722 	(WX2848,WX2845,WX2846);
	or 	XG16723 	(WX2862,WX2859,WX2860);
	or 	XG16724 	(WX2876,WX2873,WX2874);
	or 	XG16725 	(WX2890,WX2887,WX2888);
	or 	XG16726 	(WX2904,WX2901,WX2902);
	or 	XG16727 	(WX2918,WX2915,WX2916);
	or 	XG16728 	(WX2932,WX2929,WX2930);
	or 	XG16729 	(WX2946,WX2943,WX2944);
	or 	XG16730 	(WX2960,WX2957,WX2958);
	or 	XG16731 	(WX2974,WX2971,WX2972);
	or 	XG16732 	(WX2988,WX2985,WX2986);
	or 	XG16733 	(WX3002,WX2999,WX3000);
	or 	XG16734 	(WX3016,WX3013,WX3014);
	or 	XG16735 	(WX3030,WX3027,WX3028);
	or 	XG16736 	(WX3044,WX3041,WX3042);
	or 	XG16737 	(WX3058,WX3055,WX3056);
	or 	XG16738 	(WX3917,WX3914,WX3915);
	or 	XG16739 	(WX3931,WX3928,WX3929);
	or 	XG16740 	(WX3945,WX3942,WX3943);
	or 	XG16741 	(WX3959,WX3956,WX3957);
	or 	XG16742 	(WX3973,WX3970,WX3971);
	or 	XG16743 	(WX3987,WX3984,WX3985);
	or 	XG16744 	(WX4001,WX3998,WX3999);
	or 	XG16745 	(WX4015,WX4012,WX4013);
	or 	XG16746 	(WX4029,WX4026,WX4027);
	or 	XG16747 	(WX4043,WX4040,WX4041);
	or 	XG16748 	(WX4057,WX4054,WX4055);
	or 	XG16749 	(WX4071,WX4068,WX4069);
	or 	XG16750 	(WX4085,WX4082,WX4083);
	or 	XG16751 	(WX4099,WX4096,WX4097);
	or 	XG16752 	(WX4113,WX4110,WX4111);
	or 	XG16753 	(WX4127,WX4124,WX4125);
	or 	XG16754 	(WX4141,WX4138,WX4139);
	or 	XG16755 	(WX4155,WX4152,WX4153);
	or 	XG16756 	(WX4169,WX4166,WX4167);
	or 	XG16757 	(WX4183,WX4180,WX4181);
	or 	XG16758 	(WX4197,WX4194,WX4195);
	or 	XG16759 	(WX4211,WX4208,WX4209);
	or 	XG16760 	(WX4225,WX4222,WX4223);
	or 	XG16761 	(WX4239,WX4236,WX4237);
	or 	XG16762 	(WX4253,WX4250,WX4251);
	or 	XG16763 	(WX4267,WX4264,WX4265);
	or 	XG16764 	(WX4281,WX4278,WX4279);
	or 	XG16765 	(WX4295,WX4292,WX4293);
	or 	XG16766 	(WX4309,WX4306,WX4307);
	or 	XG16767 	(WX4323,WX4320,WX4321);
	or 	XG16768 	(WX4337,WX4334,WX4335);
	or 	XG16769 	(WX4351,WX4348,WX4349);
	or 	XG16770 	(WX5210,WX5207,WX5208);
	or 	XG16771 	(WX5224,WX5221,WX5222);
	or 	XG16772 	(WX5238,WX5235,WX5236);
	or 	XG16773 	(WX5252,WX5249,WX5250);
	or 	XG16774 	(WX5266,WX5263,WX5264);
	or 	XG16775 	(WX5280,WX5277,WX5278);
	or 	XG16776 	(WX5294,WX5291,WX5292);
	or 	XG16777 	(WX5308,WX5305,WX5306);
	or 	XG16778 	(WX5322,WX5319,WX5320);
	or 	XG16779 	(WX5336,WX5333,WX5334);
	or 	XG16780 	(WX5350,WX5347,WX5348);
	or 	XG16781 	(WX5364,WX5361,WX5362);
	or 	XG16782 	(WX5378,WX5375,WX5376);
	or 	XG16783 	(WX5392,WX5389,WX5390);
	or 	XG16784 	(WX5406,WX5403,WX5404);
	or 	XG16785 	(WX5420,WX5417,WX5418);
	or 	XG16786 	(WX5434,WX5431,WX5432);
	or 	XG16787 	(WX5448,WX5445,WX5446);
	or 	XG16788 	(WX5462,WX5459,WX5460);
	or 	XG16789 	(WX5476,WX5473,WX5474);
	or 	XG16790 	(WX5490,WX5487,WX5488);
	or 	XG16791 	(WX5504,WX5501,WX5502);
	or 	XG16792 	(WX5518,WX5515,WX5516);
	or 	XG16793 	(WX5532,WX5529,WX5530);
	or 	XG16794 	(WX5546,WX5543,WX5544);
	or 	XG16795 	(WX5560,WX5557,WX5558);
	or 	XG16796 	(WX5574,WX5571,WX5572);
	or 	XG16797 	(WX5588,WX5585,WX5586);
	or 	XG16798 	(WX5602,WX5599,WX5600);
	or 	XG16799 	(WX5616,WX5613,WX5614);
	or 	XG16800 	(WX5630,WX5627,WX5628);
	or 	XG16801 	(WX5644,WX5641,WX5642);
	or 	XG16802 	(WX6503,WX6500,WX6501);
	or 	XG16803 	(WX6517,WX6514,WX6515);
	or 	XG16804 	(WX6531,WX6528,WX6529);
	or 	XG16805 	(WX6545,WX6542,WX6543);
	or 	XG16806 	(WX6559,WX6556,WX6557);
	or 	XG16807 	(WX6573,WX6570,WX6571);
	or 	XG16808 	(WX6587,WX6584,WX6585);
	or 	XG16809 	(WX6601,WX6598,WX6599);
	or 	XG16810 	(WX6615,WX6612,WX6613);
	or 	XG16811 	(WX6629,WX6626,WX6627);
	or 	XG16812 	(WX6643,WX6640,WX6641);
	or 	XG16813 	(WX6657,WX6654,WX6655);
	or 	XG16814 	(WX6671,WX6668,WX6669);
	or 	XG16815 	(WX6685,WX6682,WX6683);
	or 	XG16816 	(WX6699,WX6696,WX6697);
	or 	XG16817 	(WX6713,WX6710,WX6711);
	or 	XG16818 	(WX6727,WX6724,WX6725);
	or 	XG16819 	(WX6741,WX6738,WX6739);
	or 	XG16820 	(WX6755,WX6752,WX6753);
	or 	XG16821 	(WX6769,WX6766,WX6767);
	or 	XG16822 	(WX6783,WX6780,WX6781);
	or 	XG16823 	(WX6797,WX6794,WX6795);
	or 	XG16824 	(WX6811,WX6808,WX6809);
	or 	XG16825 	(WX6825,WX6822,WX6823);
	or 	XG16826 	(WX6839,WX6836,WX6837);
	or 	XG16827 	(WX6853,WX6850,WX6851);
	or 	XG16828 	(WX6867,WX6864,WX6865);
	or 	XG16829 	(WX6881,WX6878,WX6879);
	or 	XG16830 	(WX6895,WX6892,WX6893);
	or 	XG16831 	(WX6909,WX6906,WX6907);
	or 	XG16832 	(WX6923,WX6920,WX6921);
	or 	XG16833 	(WX6937,WX6934,WX6935);
	or 	XG16834 	(WX7796,WX7793,WX7794);
	or 	XG16835 	(WX7810,WX7807,WX7808);
	or 	XG16836 	(WX7824,WX7821,WX7822);
	or 	XG16837 	(WX7838,WX7835,WX7836);
	or 	XG16838 	(WX7852,WX7849,WX7850);
	or 	XG16839 	(WX7866,WX7863,WX7864);
	or 	XG16840 	(WX7880,WX7877,WX7878);
	or 	XG16841 	(WX7894,WX7891,WX7892);
	or 	XG16842 	(WX7908,WX7905,WX7906);
	or 	XG16843 	(WX7922,WX7919,WX7920);
	or 	XG16844 	(WX7936,WX7933,WX7934);
	or 	XG16845 	(WX7950,WX7947,WX7948);
	or 	XG16846 	(WX7964,WX7961,WX7962);
	or 	XG16847 	(WX7978,WX7975,WX7976);
	or 	XG16848 	(WX7992,WX7989,WX7990);
	or 	XG16849 	(WX8006,WX8003,WX8004);
	or 	XG16850 	(WX8020,WX8017,WX8018);
	or 	XG16851 	(WX8034,WX8031,WX8032);
	or 	XG16852 	(WX8048,WX8045,WX8046);
	or 	XG16853 	(WX8062,WX8059,WX8060);
	or 	XG16854 	(WX8076,WX8073,WX8074);
	or 	XG16855 	(WX8090,WX8087,WX8088);
	or 	XG16856 	(WX8104,WX8101,WX8102);
	or 	XG16857 	(WX8118,WX8115,WX8116);
	or 	XG16858 	(WX8132,WX8129,WX8130);
	or 	XG16859 	(WX8146,WX8143,WX8144);
	or 	XG16860 	(WX8160,WX8157,WX8158);
	or 	XG16861 	(WX8174,WX8171,WX8172);
	or 	XG16862 	(WX8188,WX8185,WX8186);
	or 	XG16863 	(WX8202,WX8199,WX8200);
	or 	XG16864 	(WX8216,WX8213,WX8214);
	or 	XG16865 	(WX8230,WX8227,WX8228);
	or 	XG16866 	(WX9089,WX9086,WX9087);
	or 	XG16867 	(WX9103,WX9100,WX9101);
	or 	XG16868 	(WX9117,WX9114,WX9115);
	or 	XG16869 	(WX9131,WX9128,WX9129);
	or 	XG16870 	(WX9145,WX9142,WX9143);
	or 	XG16871 	(WX9159,WX9156,WX9157);
	or 	XG16872 	(WX9173,WX9170,WX9171);
	or 	XG16873 	(WX9187,WX9184,WX9185);
	or 	XG16874 	(WX9201,WX9198,WX9199);
	or 	XG16875 	(WX9215,WX9212,WX9213);
	or 	XG16876 	(WX9229,WX9226,WX9227);
	or 	XG16877 	(WX9243,WX9240,WX9241);
	or 	XG16878 	(WX9257,WX9254,WX9255);
	or 	XG16879 	(WX9271,WX9268,WX9269);
	or 	XG16880 	(WX9285,WX9282,WX9283);
	or 	XG16881 	(WX9299,WX9296,WX9297);
	or 	XG16882 	(WX9313,WX9310,WX9311);
	or 	XG16883 	(WX9327,WX9324,WX9325);
	or 	XG16884 	(WX9341,WX9338,WX9339);
	or 	XG16885 	(WX9355,WX9352,WX9353);
	or 	XG16886 	(WX9369,WX9366,WX9367);
	or 	XG16887 	(WX9383,WX9380,WX9381);
	or 	XG16888 	(WX9397,WX9394,WX9395);
	or 	XG16889 	(WX9411,WX9408,WX9409);
	or 	XG16890 	(WX9425,WX9422,WX9423);
	or 	XG16891 	(WX9439,WX9436,WX9437);
	or 	XG16892 	(WX9453,WX9450,WX9451);
	or 	XG16893 	(WX9467,WX9464,WX9465);
	or 	XG16894 	(WX9481,WX9478,WX9479);
	or 	XG16895 	(WX9495,WX9492,WX9493);
	or 	XG16896 	(WX9509,WX9506,WX9507);
	or 	XG16897 	(WX9523,WX9520,WX9521);
	or 	XG16898 	(WX10382,WX10379,WX10380);
	or 	XG16899 	(WX10396,WX10393,WX10394);
	or 	XG16900 	(WX10410,WX10407,WX10408);
	or 	XG16901 	(WX10424,WX10421,WX10422);
	or 	XG16902 	(WX10438,WX10435,WX10436);
	or 	XG16903 	(WX10452,WX10449,WX10450);
	or 	XG16904 	(WX10466,WX10463,WX10464);
	or 	XG16905 	(WX10480,WX10477,WX10478);
	or 	XG16906 	(WX10494,WX10491,WX10492);
	or 	XG16907 	(WX10508,WX10505,WX10506);
	or 	XG16908 	(WX10522,WX10519,WX10520);
	or 	XG16909 	(WX10536,WX10533,WX10534);
	or 	XG16910 	(WX10550,WX10547,WX10548);
	or 	XG16911 	(WX10564,WX10561,WX10562);
	or 	XG16912 	(WX10578,WX10575,WX10576);
	or 	XG16913 	(WX10592,WX10589,WX10590);
	or 	XG16914 	(WX10606,WX10603,WX10604);
	or 	XG16915 	(WX10620,WX10617,WX10618);
	or 	XG16916 	(WX10634,WX10631,WX10632);
	or 	XG16917 	(WX10648,WX10645,WX10646);
	or 	XG16918 	(WX10662,WX10659,WX10660);
	or 	XG16919 	(WX10676,WX10673,WX10674);
	or 	XG16920 	(WX10690,WX10687,WX10688);
	or 	XG16921 	(WX10704,WX10701,WX10702);
	or 	XG16922 	(WX10718,WX10715,WX10716);
	or 	XG16923 	(WX10732,WX10729,WX10730);
	or 	XG16924 	(WX10746,WX10743,WX10744);
	or 	XG16925 	(WX10760,WX10757,WX10758);
	or 	XG16926 	(WX10774,WX10771,WX10772);
	or 	XG16927 	(WX10788,WX10785,WX10786);
	or 	XG16928 	(WX10802,WX10799,WX10800);
	or 	XG16929 	(WX10816,WX10813,WX10814);
	not 	XG16930 	(WX10825,WX10816);
	not 	XG16931 	(WX10811,WX10802);
	not 	XG16932 	(WX10797,WX10788);
	not 	XG16933 	(WX10783,WX10774);
	not 	XG16934 	(WX10769,WX10760);
	not 	XG16935 	(WX10755,WX10746);
	not 	XG16936 	(WX10741,WX10732);
	not 	XG16937 	(WX10727,WX10718);
	not 	XG16938 	(WX10713,WX10704);
	not 	XG16939 	(WX10699,WX10690);
	not 	XG16940 	(WX10685,WX10676);
	not 	XG16941 	(WX10671,WX10662);
	not 	XG16942 	(WX10657,WX10648);
	not 	XG16943 	(WX10643,WX10634);
	not 	XG16944 	(WX10629,WX10620);
	not 	XG16945 	(WX10615,WX10606);
	not 	XG16946 	(WX10601,WX10592);
	not 	XG16947 	(WX10587,WX10578);
	not 	XG16948 	(WX10573,WX10564);
	not 	XG16949 	(WX10559,WX10550);
	not 	XG16950 	(WX10545,WX10536);
	not 	XG16951 	(WX10531,WX10522);
	not 	XG16952 	(WX10517,WX10508);
	not 	XG16953 	(WX10503,WX10494);
	not 	XG16954 	(WX10489,WX10480);
	not 	XG16955 	(WX10475,WX10466);
	not 	XG16956 	(WX10461,WX10452);
	not 	XG16957 	(WX10447,WX10438);
	not 	XG16958 	(WX10433,WX10424);
	not 	XG16959 	(WX10419,WX10410);
	not 	XG16960 	(WX10405,WX10396);
	not 	XG16961 	(WX10391,WX10382);
	not 	XG16962 	(WX9532,WX9523);
	not 	XG16963 	(WX9518,WX9509);
	not 	XG16964 	(WX9504,WX9495);
	not 	XG16965 	(WX9490,WX9481);
	not 	XG16966 	(WX9476,WX9467);
	not 	XG16967 	(WX9462,WX9453);
	not 	XG16968 	(WX9448,WX9439);
	not 	XG16969 	(WX9434,WX9425);
	not 	XG16970 	(WX9420,WX9411);
	not 	XG16971 	(WX9406,WX9397);
	not 	XG16972 	(WX9392,WX9383);
	not 	XG16973 	(WX9378,WX9369);
	not 	XG16974 	(WX9364,WX9355);
	not 	XG16975 	(WX9350,WX9341);
	not 	XG16976 	(WX9336,WX9327);
	not 	XG16977 	(WX9322,WX9313);
	not 	XG16978 	(WX9308,WX9299);
	not 	XG16979 	(WX9294,WX9285);
	not 	XG16980 	(WX9280,WX9271);
	not 	XG16981 	(WX9266,WX9257);
	not 	XG16982 	(WX9252,WX9243);
	not 	XG16983 	(WX9238,WX9229);
	not 	XG16984 	(WX9224,WX9215);
	not 	XG16985 	(WX9210,WX9201);
	not 	XG16986 	(WX9196,WX9187);
	not 	XG16987 	(WX9182,WX9173);
	not 	XG16988 	(WX9168,WX9159);
	not 	XG16989 	(WX9154,WX9145);
	not 	XG16990 	(WX9140,WX9131);
	not 	XG16991 	(WX9126,WX9117);
	not 	XG16992 	(WX9112,WX9103);
	not 	XG16993 	(WX9098,WX9089);
	not 	XG16994 	(WX8239,WX8230);
	not 	XG16995 	(WX8225,WX8216);
	not 	XG16996 	(WX8211,WX8202);
	not 	XG16997 	(WX8197,WX8188);
	not 	XG16998 	(WX8183,WX8174);
	not 	XG16999 	(WX8169,WX8160);
	not 	XG17000 	(WX8155,WX8146);
	not 	XG17001 	(WX8141,WX8132);
	not 	XG17002 	(WX8127,WX8118);
	not 	XG17003 	(WX8113,WX8104);
	not 	XG17004 	(WX8099,WX8090);
	not 	XG17005 	(WX8085,WX8076);
	not 	XG17006 	(WX8071,WX8062);
	not 	XG17007 	(WX8057,WX8048);
	not 	XG17008 	(WX8043,WX8034);
	not 	XG17009 	(WX8029,WX8020);
	not 	XG17010 	(WX8015,WX8006);
	not 	XG17011 	(WX8001,WX7992);
	not 	XG17012 	(WX7987,WX7978);
	not 	XG17013 	(WX7973,WX7964);
	not 	XG17014 	(WX7959,WX7950);
	not 	XG17015 	(WX7945,WX7936);
	not 	XG17016 	(WX7931,WX7922);
	not 	XG17017 	(WX7917,WX7908);
	not 	XG17018 	(WX7903,WX7894);
	not 	XG17019 	(WX7889,WX7880);
	not 	XG17020 	(WX7875,WX7866);
	not 	XG17021 	(WX7861,WX7852);
	not 	XG17022 	(WX7847,WX7838);
	not 	XG17023 	(WX7833,WX7824);
	not 	XG17024 	(WX7819,WX7810);
	not 	XG17025 	(WX7805,WX7796);
	not 	XG17026 	(WX6946,WX6937);
	not 	XG17027 	(WX6932,WX6923);
	not 	XG17028 	(WX6918,WX6909);
	not 	XG17029 	(WX6904,WX6895);
	not 	XG17030 	(WX6890,WX6881);
	not 	XG17031 	(WX6876,WX6867);
	not 	XG17032 	(WX6862,WX6853);
	not 	XG17033 	(WX6848,WX6839);
	not 	XG17034 	(WX6834,WX6825);
	not 	XG17035 	(WX6820,WX6811);
	not 	XG17036 	(WX6806,WX6797);
	not 	XG17037 	(WX6792,WX6783);
	not 	XG17038 	(WX6778,WX6769);
	not 	XG17039 	(WX6764,WX6755);
	not 	XG17040 	(WX6750,WX6741);
	not 	XG17041 	(WX6736,WX6727);
	not 	XG17042 	(WX6722,WX6713);
	not 	XG17043 	(WX6708,WX6699);
	not 	XG17044 	(WX6694,WX6685);
	not 	XG17045 	(WX6680,WX6671);
	not 	XG17046 	(WX6666,WX6657);
	not 	XG17047 	(WX6652,WX6643);
	not 	XG17048 	(WX6638,WX6629);
	not 	XG17049 	(WX6624,WX6615);
	not 	XG17050 	(WX6610,WX6601);
	not 	XG17051 	(WX6596,WX6587);
	not 	XG17052 	(WX6582,WX6573);
	not 	XG17053 	(WX6568,WX6559);
	not 	XG17054 	(WX6554,WX6545);
	not 	XG17055 	(WX6540,WX6531);
	not 	XG17056 	(WX6526,WX6517);
	not 	XG17057 	(WX6512,WX6503);
	not 	XG17058 	(WX5653,WX5644);
	not 	XG17059 	(WX5639,WX5630);
	not 	XG17060 	(WX5625,WX5616);
	not 	XG17061 	(WX5611,WX5602);
	not 	XG17062 	(WX5597,WX5588);
	not 	XG17063 	(WX5583,WX5574);
	not 	XG17064 	(WX5569,WX5560);
	not 	XG17065 	(WX5555,WX5546);
	not 	XG17066 	(WX5541,WX5532);
	not 	XG17067 	(WX5527,WX5518);
	not 	XG17068 	(WX5513,WX5504);
	not 	XG17069 	(WX5499,WX5490);
	not 	XG17070 	(WX5485,WX5476);
	not 	XG17071 	(WX5471,WX5462);
	not 	XG17072 	(WX5457,WX5448);
	not 	XG17073 	(WX5443,WX5434);
	not 	XG17074 	(WX5429,WX5420);
	not 	XG17075 	(WX5415,WX5406);
	not 	XG17076 	(WX5401,WX5392);
	not 	XG17077 	(WX5387,WX5378);
	not 	XG17078 	(WX5373,WX5364);
	not 	XG17079 	(WX5359,WX5350);
	not 	XG17080 	(WX5345,WX5336);
	not 	XG17081 	(WX5331,WX5322);
	not 	XG17082 	(WX5317,WX5308);
	not 	XG17083 	(WX5303,WX5294);
	not 	XG17084 	(WX5289,WX5280);
	not 	XG17085 	(WX5275,WX5266);
	not 	XG17086 	(WX5261,WX5252);
	not 	XG17087 	(WX5247,WX5238);
	not 	XG17088 	(WX5233,WX5224);
	not 	XG17089 	(WX5219,WX5210);
	not 	XG17090 	(WX4360,WX4351);
	not 	XG17091 	(WX4346,WX4337);
	not 	XG17092 	(WX4332,WX4323);
	not 	XG17093 	(WX4318,WX4309);
	not 	XG17094 	(WX4304,WX4295);
	not 	XG17095 	(WX4290,WX4281);
	not 	XG17096 	(WX4276,WX4267);
	not 	XG17097 	(WX4262,WX4253);
	not 	XG17098 	(WX4248,WX4239);
	not 	XG17099 	(WX4234,WX4225);
	not 	XG17100 	(WX4220,WX4211);
	not 	XG17101 	(WX4206,WX4197);
	not 	XG17102 	(WX4192,WX4183);
	not 	XG17103 	(WX4178,WX4169);
	not 	XG17104 	(WX4164,WX4155);
	not 	XG17105 	(WX4150,WX4141);
	not 	XG17106 	(WX4136,WX4127);
	not 	XG17107 	(WX4122,WX4113);
	not 	XG17108 	(WX4108,WX4099);
	not 	XG17109 	(WX4094,WX4085);
	not 	XG17110 	(WX4080,WX4071);
	not 	XG17111 	(WX4066,WX4057);
	not 	XG17112 	(WX4052,WX4043);
	not 	XG17113 	(WX4038,WX4029);
	not 	XG17114 	(WX4024,WX4015);
	not 	XG17115 	(WX4010,WX4001);
	not 	XG17116 	(WX3996,WX3987);
	not 	XG17117 	(WX3982,WX3973);
	not 	XG17118 	(WX3968,WX3959);
	not 	XG17119 	(WX3954,WX3945);
	not 	XG17120 	(WX3940,WX3931);
	not 	XG17121 	(WX3926,WX3917);
	not 	XG17122 	(WX3067,WX3058);
	not 	XG17123 	(WX3053,WX3044);
	not 	XG17124 	(WX3039,WX3030);
	not 	XG17125 	(WX3025,WX3016);
	not 	XG17126 	(WX3011,WX3002);
	not 	XG17127 	(WX2997,WX2988);
	not 	XG17128 	(WX2983,WX2974);
	not 	XG17129 	(WX2969,WX2960);
	not 	XG17130 	(WX2955,WX2946);
	not 	XG17131 	(WX2941,WX2932);
	not 	XG17132 	(WX2927,WX2918);
	not 	XG17133 	(WX2913,WX2904);
	not 	XG17134 	(WX2899,WX2890);
	not 	XG17135 	(WX2885,WX2876);
	not 	XG17136 	(WX2871,WX2862);
	not 	XG17137 	(WX2857,WX2848);
	not 	XG17138 	(WX2843,WX2834);
	not 	XG17139 	(WX2829,WX2820);
	not 	XG17140 	(WX2815,WX2806);
	not 	XG17141 	(WX2801,WX2792);
	not 	XG17142 	(WX2787,WX2778);
	not 	XG17143 	(WX2773,WX2764);
	not 	XG17144 	(WX2759,WX2750);
	not 	XG17145 	(WX2745,WX2736);
	not 	XG17146 	(WX2731,WX2722);
	not 	XG17147 	(WX2717,WX2708);
	not 	XG17148 	(WX2703,WX2694);
	not 	XG17149 	(WX2689,WX2680);
	not 	XG17150 	(WX2675,WX2666);
	not 	XG17151 	(WX2661,WX2652);
	not 	XG17152 	(WX2647,WX2638);
	not 	XG17153 	(WX2633,WX2624);
	not 	XG17154 	(WX1774,WX1765);
	not 	XG17155 	(WX1760,WX1751);
	not 	XG17156 	(WX1746,WX1737);
	not 	XG17157 	(WX1732,WX1723);
	not 	XG17158 	(WX1718,WX1709);
	not 	XG17159 	(WX1704,WX1695);
	not 	XG17160 	(WX1690,WX1681);
	not 	XG17161 	(WX1676,WX1667);
	not 	XG17162 	(WX1662,WX1653);
	not 	XG17163 	(WX1648,WX1639);
	not 	XG17164 	(WX1634,WX1625);
	not 	XG17165 	(WX1620,WX1611);
	not 	XG17166 	(WX1606,WX1597);
	not 	XG17167 	(WX1592,WX1583);
	not 	XG17168 	(WX1578,WX1569);
	not 	XG17169 	(WX1564,WX1555);
	not 	XG17170 	(WX1550,WX1541);
	not 	XG17171 	(WX1536,WX1527);
	not 	XG17172 	(WX1522,WX1513);
	not 	XG17173 	(WX1508,WX1499);
	not 	XG17174 	(WX1494,WX1485);
	not 	XG17175 	(WX1480,WX1471);
	not 	XG17176 	(WX1466,WX1457);
	not 	XG17177 	(WX1452,WX1443);
	not 	XG17178 	(WX1438,WX1429);
	not 	XG17179 	(WX1424,WX1415);
	not 	XG17180 	(WX1410,WX1401);
	not 	XG17181 	(WX1396,WX1387);
	not 	XG17182 	(WX1382,WX1373);
	not 	XG17183 	(WX1368,WX1359);
	not 	XG17184 	(WX1354,WX1345);
	not 	XG17185 	(WX1340,WX1331);
	not 	XG17186 	(WX481,WX472);
	not 	XG17187 	(WX467,WX458);
	not 	XG17188 	(WX453,WX444);
	not 	XG17189 	(WX439,WX430);
	not 	XG17190 	(WX425,WX416);
	not 	XG17191 	(WX411,WX402);
	not 	XG17192 	(WX397,WX388);
	not 	XG17193 	(WX383,WX374);
	not 	XG17194 	(WX369,WX360);
	not 	XG17195 	(WX355,WX346);
	not 	XG17196 	(WX341,WX332);
	not 	XG17197 	(WX327,WX318);
	not 	XG17198 	(WX313,WX304);
	not 	XG17199 	(WX299,WX290);
	not 	XG17200 	(WX285,WX276);
	not 	XG17201 	(WX271,WX262);
	not 	XG17202 	(WX257,WX248);
	not 	XG17203 	(WX243,WX234);
	not 	XG17204 	(WX229,WX220);
	not 	XG17205 	(WX215,WX206);
	not 	XG17206 	(WX201,WX192);
	not 	XG17207 	(WX187,WX178);
	not 	XG17208 	(WX173,WX164);
	not 	XG17209 	(WX159,WX150);
	not 	XG17210 	(WX145,WX136);
	not 	XG17211 	(WX131,WX122);
	not 	XG17212 	(WX117,WX108);
	not 	XG17213 	(WX103,WX94);
	not 	XG17214 	(WX89,WX80);
	not 	XG17215 	(WX75,WX66);
	not 	XG17216 	(WX61,WX52);
	not 	XG17217 	(WX47,WX38);
	not 	XG17218 	(WX48,WX47);
	not 	XG17219 	(WX62,WX61);
	not 	XG17220 	(WX76,WX75);
	not 	XG17221 	(WX90,WX89);
	not 	XG17222 	(WX104,WX103);
	not 	XG17223 	(WX118,WX117);
	not 	XG17224 	(WX132,WX131);
	not 	XG17225 	(WX146,WX145);
	not 	XG17226 	(WX160,WX159);
	not 	XG17227 	(WX174,WX173);
	not 	XG17228 	(WX188,WX187);
	not 	XG17229 	(WX202,WX201);
	not 	XG17230 	(WX216,WX215);
	not 	XG17231 	(WX230,WX229);
	not 	XG17232 	(WX244,WX243);
	not 	XG17233 	(WX258,WX257);
	not 	XG17234 	(WX272,WX271);
	not 	XG17235 	(WX286,WX285);
	not 	XG17236 	(WX300,WX299);
	not 	XG17237 	(WX314,WX313);
	not 	XG17238 	(WX328,WX327);
	not 	XG17239 	(WX342,WX341);
	not 	XG17240 	(WX356,WX355);
	not 	XG17241 	(WX370,WX369);
	not 	XG17242 	(WX384,WX383);
	not 	XG17243 	(WX398,WX397);
	not 	XG17244 	(WX412,WX411);
	not 	XG17245 	(WX426,WX425);
	not 	XG17246 	(WX440,WX439);
	not 	XG17247 	(WX454,WX453);
	not 	XG17248 	(WX468,WX467);
	not 	XG17249 	(WX482,WX481);
	not 	XG17250 	(WX1341,WX1340);
	not 	XG17251 	(WX1355,WX1354);
	not 	XG17252 	(WX1369,WX1368);
	not 	XG17253 	(WX1383,WX1382);
	not 	XG17254 	(WX1397,WX1396);
	not 	XG17255 	(WX1411,WX1410);
	not 	XG17256 	(WX1425,WX1424);
	not 	XG17257 	(WX1439,WX1438);
	not 	XG17258 	(WX1453,WX1452);
	not 	XG17259 	(WX1467,WX1466);
	not 	XG17260 	(WX1481,WX1480);
	not 	XG17261 	(WX1495,WX1494);
	not 	XG17262 	(WX1509,WX1508);
	not 	XG17263 	(WX1523,WX1522);
	not 	XG17264 	(WX1537,WX1536);
	not 	XG17265 	(WX1551,WX1550);
	not 	XG17266 	(WX1565,WX1564);
	not 	XG17267 	(WX1579,WX1578);
	not 	XG17268 	(WX1593,WX1592);
	not 	XG17269 	(WX1607,WX1606);
	not 	XG17270 	(WX1621,WX1620);
	not 	XG17271 	(WX1635,WX1634);
	not 	XG17272 	(WX1649,WX1648);
	not 	XG17273 	(WX1663,WX1662);
	not 	XG17274 	(WX1677,WX1676);
	not 	XG17275 	(WX1691,WX1690);
	not 	XG17276 	(WX1705,WX1704);
	not 	XG17277 	(WX1719,WX1718);
	not 	XG17278 	(WX1733,WX1732);
	not 	XG17279 	(WX1747,WX1746);
	not 	XG17280 	(WX1761,WX1760);
	not 	XG17281 	(WX1775,WX1774);
	not 	XG17282 	(WX2634,WX2633);
	not 	XG17283 	(WX2648,WX2647);
	not 	XG17284 	(WX2662,WX2661);
	not 	XG17285 	(WX2676,WX2675);
	not 	XG17286 	(WX2690,WX2689);
	not 	XG17287 	(WX2704,WX2703);
	not 	XG17288 	(WX2718,WX2717);
	not 	XG17289 	(WX2732,WX2731);
	not 	XG17290 	(WX2746,WX2745);
	not 	XG17291 	(WX2760,WX2759);
	not 	XG17292 	(WX2774,WX2773);
	not 	XG17293 	(WX2788,WX2787);
	not 	XG17294 	(WX2802,WX2801);
	not 	XG17295 	(WX2816,WX2815);
	not 	XG17296 	(WX2830,WX2829);
	not 	XG17297 	(WX2844,WX2843);
	not 	XG17298 	(WX2858,WX2857);
	not 	XG17299 	(WX2872,WX2871);
	not 	XG17300 	(WX2886,WX2885);
	not 	XG17301 	(WX2900,WX2899);
	not 	XG17302 	(WX2914,WX2913);
	not 	XG17303 	(WX2928,WX2927);
	not 	XG17304 	(WX2942,WX2941);
	not 	XG17305 	(WX2956,WX2955);
	not 	XG17306 	(WX2970,WX2969);
	not 	XG17307 	(WX2984,WX2983);
	not 	XG17308 	(WX2998,WX2997);
	not 	XG17309 	(WX3012,WX3011);
	not 	XG17310 	(WX3026,WX3025);
	not 	XG17311 	(WX3040,WX3039);
	not 	XG17312 	(WX3054,WX3053);
	not 	XG17313 	(WX3068,WX3067);
	not 	XG17314 	(WX3927,WX3926);
	not 	XG17315 	(WX3941,WX3940);
	not 	XG17316 	(WX3955,WX3954);
	not 	XG17317 	(WX3969,WX3968);
	not 	XG17318 	(WX3983,WX3982);
	not 	XG17319 	(WX3997,WX3996);
	not 	XG17320 	(WX4011,WX4010);
	not 	XG17321 	(WX4025,WX4024);
	not 	XG17322 	(WX4039,WX4038);
	not 	XG17323 	(WX4053,WX4052);
	not 	XG17324 	(WX4067,WX4066);
	not 	XG17325 	(WX4081,WX4080);
	not 	XG17326 	(WX4095,WX4094);
	not 	XG17327 	(WX4109,WX4108);
	not 	XG17328 	(WX4123,WX4122);
	not 	XG17329 	(WX4137,WX4136);
	not 	XG17330 	(WX4151,WX4150);
	not 	XG17331 	(WX4165,WX4164);
	not 	XG17332 	(WX4179,WX4178);
	not 	XG17333 	(WX4193,WX4192);
	not 	XG17334 	(WX4207,WX4206);
	not 	XG17335 	(WX4221,WX4220);
	not 	XG17336 	(WX4235,WX4234);
	not 	XG17337 	(WX4249,WX4248);
	not 	XG17338 	(WX4263,WX4262);
	not 	XG17339 	(WX4277,WX4276);
	not 	XG17340 	(WX4291,WX4290);
	not 	XG17341 	(WX4305,WX4304);
	not 	XG17342 	(WX4319,WX4318);
	not 	XG17343 	(WX4333,WX4332);
	not 	XG17344 	(WX4347,WX4346);
	not 	XG17345 	(WX4361,WX4360);
	not 	XG17346 	(WX5220,WX5219);
	not 	XG17347 	(WX5234,WX5233);
	not 	XG17348 	(WX5248,WX5247);
	not 	XG17349 	(WX5262,WX5261);
	not 	XG17350 	(WX5276,WX5275);
	not 	XG17351 	(WX5290,WX5289);
	not 	XG17352 	(WX5304,WX5303);
	not 	XG17353 	(WX5318,WX5317);
	not 	XG17354 	(WX5332,WX5331);
	not 	XG17355 	(WX5346,WX5345);
	not 	XG17356 	(WX5360,WX5359);
	not 	XG17357 	(WX5374,WX5373);
	not 	XG17358 	(WX5388,WX5387);
	not 	XG17359 	(WX5402,WX5401);
	not 	XG17360 	(WX5416,WX5415);
	not 	XG17361 	(WX5430,WX5429);
	not 	XG17362 	(WX5444,WX5443);
	not 	XG17363 	(WX5458,WX5457);
	not 	XG17364 	(WX5472,WX5471);
	not 	XG17365 	(WX5486,WX5485);
	not 	XG17366 	(WX5500,WX5499);
	not 	XG17367 	(WX5514,WX5513);
	not 	XG17368 	(WX5528,WX5527);
	not 	XG17369 	(WX5542,WX5541);
	not 	XG17370 	(WX5556,WX5555);
	not 	XG17371 	(WX5570,WX5569);
	not 	XG17372 	(WX5584,WX5583);
	not 	XG17373 	(WX5598,WX5597);
	not 	XG17374 	(WX5612,WX5611);
	not 	XG17375 	(WX5626,WX5625);
	not 	XG17376 	(WX5640,WX5639);
	not 	XG17377 	(WX5654,WX5653);
	not 	XG17378 	(WX6513,WX6512);
	not 	XG17379 	(WX6527,WX6526);
	not 	XG17380 	(WX6541,WX6540);
	not 	XG17381 	(WX6555,WX6554);
	not 	XG17382 	(WX6569,WX6568);
	not 	XG17383 	(WX6583,WX6582);
	not 	XG17384 	(WX6597,WX6596);
	not 	XG17385 	(WX6611,WX6610);
	not 	XG17386 	(WX6625,WX6624);
	not 	XG17387 	(WX6639,WX6638);
	not 	XG17388 	(WX6653,WX6652);
	not 	XG17389 	(WX6667,WX6666);
	not 	XG17390 	(WX6681,WX6680);
	not 	XG17391 	(WX6695,WX6694);
	not 	XG17392 	(WX6709,WX6708);
	not 	XG17393 	(WX6723,WX6722);
	not 	XG17394 	(WX6737,WX6736);
	not 	XG17395 	(WX6751,WX6750);
	not 	XG17396 	(WX6765,WX6764);
	not 	XG17397 	(WX6779,WX6778);
	not 	XG17398 	(WX6793,WX6792);
	not 	XG17399 	(WX6807,WX6806);
	not 	XG17400 	(WX6821,WX6820);
	not 	XG17401 	(WX6835,WX6834);
	not 	XG17402 	(WX6849,WX6848);
	not 	XG17403 	(WX6863,WX6862);
	not 	XG17404 	(WX6877,WX6876);
	not 	XG17405 	(WX6891,WX6890);
	not 	XG17406 	(WX6905,WX6904);
	not 	XG17407 	(WX6919,WX6918);
	not 	XG17408 	(WX6933,WX6932);
	not 	XG17409 	(WX6947,WX6946);
	not 	XG17410 	(WX7806,WX7805);
	not 	XG17411 	(WX7820,WX7819);
	not 	XG17412 	(WX7834,WX7833);
	not 	XG17413 	(WX7848,WX7847);
	not 	XG17414 	(WX7862,WX7861);
	not 	XG17415 	(WX7876,WX7875);
	not 	XG17416 	(WX7890,WX7889);
	not 	XG17417 	(WX7904,WX7903);
	not 	XG17418 	(WX7918,WX7917);
	not 	XG17419 	(WX7932,WX7931);
	not 	XG17420 	(WX7946,WX7945);
	not 	XG17421 	(WX7960,WX7959);
	not 	XG17422 	(WX7974,WX7973);
	not 	XG17423 	(WX7988,WX7987);
	not 	XG17424 	(WX8002,WX8001);
	not 	XG17425 	(WX8016,WX8015);
	not 	XG17426 	(WX8030,WX8029);
	not 	XG17427 	(WX8044,WX8043);
	not 	XG17428 	(WX8058,WX8057);
	not 	XG17429 	(WX8072,WX8071);
	not 	XG17430 	(WX8086,WX8085);
	not 	XG17431 	(WX8100,WX8099);
	not 	XG17432 	(WX8114,WX8113);
	not 	XG17433 	(WX8128,WX8127);
	not 	XG17434 	(WX8142,WX8141);
	not 	XG17435 	(WX8156,WX8155);
	not 	XG17436 	(WX8170,WX8169);
	not 	XG17437 	(WX8184,WX8183);
	not 	XG17438 	(WX8198,WX8197);
	not 	XG17439 	(WX8212,WX8211);
	not 	XG17440 	(WX8226,WX8225);
	not 	XG17441 	(WX8240,WX8239);
	not 	XG17442 	(WX9099,WX9098);
	not 	XG17443 	(WX9113,WX9112);
	not 	XG17444 	(WX9127,WX9126);
	not 	XG17445 	(WX9141,WX9140);
	not 	XG17446 	(WX9155,WX9154);
	not 	XG17447 	(WX9169,WX9168);
	not 	XG17448 	(WX9183,WX9182);
	not 	XG17449 	(WX9197,WX9196);
	not 	XG17450 	(WX9211,WX9210);
	not 	XG17451 	(WX9225,WX9224);
	not 	XG17452 	(WX9239,WX9238);
	not 	XG17453 	(WX9253,WX9252);
	not 	XG17454 	(WX9267,WX9266);
	not 	XG17455 	(WX9281,WX9280);
	not 	XG17456 	(WX9295,WX9294);
	not 	XG17457 	(WX9309,WX9308);
	not 	XG17458 	(WX9323,WX9322);
	not 	XG17459 	(WX9337,WX9336);
	not 	XG17460 	(WX9351,WX9350);
	not 	XG17461 	(WX9365,WX9364);
	not 	XG17462 	(WX9379,WX9378);
	not 	XG17463 	(WX9393,WX9392);
	not 	XG17464 	(WX9407,WX9406);
	not 	XG17465 	(WX9421,WX9420);
	not 	XG17466 	(WX9435,WX9434);
	not 	XG17467 	(WX9449,WX9448);
	not 	XG17468 	(WX9463,WX9462);
	not 	XG17469 	(WX9477,WX9476);
	not 	XG17470 	(WX9491,WX9490);
	not 	XG17471 	(WX9505,WX9504);
	not 	XG17472 	(WX9519,WX9518);
	not 	XG17473 	(WX9533,WX9532);
	not 	XG17474 	(WX10392,WX10391);
	not 	XG17475 	(WX10406,WX10405);
	not 	XG17476 	(WX10420,WX10419);
	not 	XG17477 	(WX10434,WX10433);
	not 	XG17478 	(WX10448,WX10447);
	not 	XG17479 	(WX10462,WX10461);
	not 	XG17480 	(WX10476,WX10475);
	not 	XG17481 	(WX10490,WX10489);
	not 	XG17482 	(WX10504,WX10503);
	not 	XG17483 	(WX10518,WX10517);
	not 	XG17484 	(WX10532,WX10531);
	not 	XG17485 	(WX10546,WX10545);
	not 	XG17486 	(WX10560,WX10559);
	not 	XG17487 	(WX10574,WX10573);
	not 	XG17488 	(WX10588,WX10587);
	not 	XG17489 	(WX10602,WX10601);
	not 	XG17490 	(WX10616,WX10615);
	not 	XG17491 	(WX10630,WX10629);
	not 	XG17492 	(WX10644,WX10643);
	not 	XG17493 	(WX10658,WX10657);
	not 	XG17494 	(WX10672,WX10671);
	not 	XG17495 	(WX10686,WX10685);
	not 	XG17496 	(WX10700,WX10699);
	not 	XG17497 	(WX10714,WX10713);
	not 	XG17498 	(WX10728,WX10727);
	not 	XG17499 	(WX10742,WX10741);
	not 	XG17500 	(WX10756,WX10755);
	not 	XG17501 	(WX10770,WX10769);
	not 	XG17502 	(WX10784,WX10783);
	not 	XG17503 	(WX10798,WX10797);
	not 	XG17504 	(WX10812,WX10811);
	not 	XG17505 	(WX10826,WX10825);
	and 	XG17506 	(WX11050,RESET,WX10826);
	and 	XG17507 	(WX11048,RESET,WX10812);
	and 	XG17508 	(WX11046,RESET,WX10798);
	and 	XG17509 	(WX11044,RESET,WX10784);
	and 	XG17510 	(WX11042,RESET,WX10770);
	and 	XG17511 	(WX11040,RESET,WX10756);
	and 	XG17512 	(WX11038,RESET,WX10742);
	and 	XG17513 	(WX11036,RESET,WX10728);
	and 	XG17514 	(WX11034,RESET,WX10714);
	and 	XG17515 	(WX11032,RESET,WX10700);
	and 	XG17516 	(WX11030,RESET,WX10686);
	and 	XG17517 	(WX11028,RESET,WX10672);
	and 	XG17518 	(WX11026,RESET,WX10658);
	and 	XG17519 	(WX11024,RESET,WX10644);
	and 	XG17520 	(WX11022,RESET,WX10630);
	and 	XG17521 	(WX11020,RESET,WX10616);
	and 	XG17522 	(WX11018,RESET,WX10602);
	and 	XG17523 	(WX11016,RESET,WX10588);
	and 	XG17524 	(WX11014,RESET,WX10574);
	and 	XG17525 	(WX11012,RESET,WX10560);
	and 	XG17526 	(WX11010,RESET,WX10546);
	and 	XG17527 	(WX11008,RESET,WX10532);
	and 	XG17528 	(WX11006,RESET,WX10518);
	and 	XG17529 	(WX11004,RESET,WX10504);
	and 	XG17530 	(WX11002,RESET,WX10490);
	and 	XG17531 	(WX11000,RESET,WX10476);
	and 	XG17532 	(WX10998,RESET,WX10462);
	and 	XG17533 	(WX10996,RESET,WX10448);
	and 	XG17534 	(WX10994,RESET,WX10434);
	and 	XG17535 	(WX10992,RESET,WX10420);
	and 	XG17536 	(WX10990,RESET,WX10406);
	and 	XG17537 	(WX10988,RESET,WX10392);
	and 	XG17538 	(WX9757,RESET,WX9533);
	and 	XG17539 	(WX9755,RESET,WX9519);
	and 	XG17540 	(WX9753,RESET,WX9505);
	and 	XG17541 	(WX9751,RESET,WX9491);
	and 	XG17542 	(WX9749,RESET,WX9477);
	and 	XG17543 	(WX9747,RESET,WX9463);
	and 	XG17544 	(WX9745,RESET,WX9449);
	and 	XG17545 	(WX9743,RESET,WX9435);
	and 	XG17546 	(WX9741,RESET,WX9421);
	and 	XG17547 	(WX9739,RESET,WX9407);
	and 	XG17548 	(WX9737,RESET,WX9393);
	and 	XG17549 	(WX9735,RESET,WX9379);
	and 	XG17550 	(WX9733,RESET,WX9365);
	and 	XG17551 	(WX9731,RESET,WX9351);
	and 	XG17552 	(WX9729,RESET,WX9337);
	and 	XG17553 	(WX9727,RESET,WX9323);
	and 	XG17554 	(WX9725,RESET,WX9309);
	and 	XG17555 	(WX9723,RESET,WX9295);
	and 	XG17556 	(WX9721,RESET,WX9281);
	and 	XG17557 	(WX9719,RESET,WX9267);
	and 	XG17558 	(WX9717,RESET,WX9253);
	and 	XG17559 	(WX9715,RESET,WX9239);
	and 	XG17560 	(WX9713,RESET,WX9225);
	and 	XG17561 	(WX9711,RESET,WX9211);
	and 	XG17562 	(WX9709,RESET,WX9197);
	and 	XG17563 	(WX9707,RESET,WX9183);
	and 	XG17564 	(WX9705,RESET,WX9169);
	and 	XG17565 	(WX9703,RESET,WX9155);
	and 	XG17566 	(WX9701,RESET,WX9141);
	and 	XG17567 	(WX9699,RESET,WX9127);
	and 	XG17568 	(WX9697,RESET,WX9113);
	and 	XG17569 	(WX9695,RESET,WX9099);
	and 	XG17570 	(WX8464,RESET,WX8240);
	and 	XG17571 	(WX8462,RESET,WX8226);
	and 	XG17572 	(WX8460,RESET,WX8212);
	and 	XG17573 	(WX8458,RESET,WX8198);
	and 	XG17574 	(WX8456,RESET,WX8184);
	and 	XG17575 	(WX8454,RESET,WX8170);
	and 	XG17576 	(WX8452,RESET,WX8156);
	and 	XG17577 	(WX8450,RESET,WX8142);
	and 	XG17578 	(WX8448,RESET,WX8128);
	and 	XG17579 	(WX8446,RESET,WX8114);
	and 	XG17580 	(WX8444,RESET,WX8100);
	and 	XG17581 	(WX8442,RESET,WX8086);
	and 	XG17582 	(WX8440,RESET,WX8072);
	and 	XG17583 	(WX8438,RESET,WX8058);
	and 	XG17584 	(WX8436,RESET,WX8044);
	and 	XG17585 	(WX8434,RESET,WX8030);
	and 	XG17586 	(WX8432,RESET,WX8016);
	and 	XG17587 	(WX8430,RESET,WX8002);
	and 	XG17588 	(WX8428,RESET,WX7988);
	and 	XG17589 	(WX8426,RESET,WX7974);
	and 	XG17590 	(WX8424,RESET,WX7960);
	and 	XG17591 	(WX8422,RESET,WX7946);
	and 	XG17592 	(WX8420,RESET,WX7932);
	and 	XG17593 	(WX8418,RESET,WX7918);
	and 	XG17594 	(WX8416,RESET,WX7904);
	and 	XG17595 	(WX8414,RESET,WX7890);
	and 	XG17596 	(WX8412,RESET,WX7876);
	and 	XG17597 	(WX8410,RESET,WX7862);
	and 	XG17598 	(WX8408,RESET,WX7848);
	and 	XG17599 	(WX8406,RESET,WX7834);
	and 	XG17600 	(WX8404,RESET,WX7820);
	and 	XG17601 	(WX8402,RESET,WX7806);
	and 	XG17602 	(WX7171,RESET,WX6947);
	and 	XG17603 	(WX7169,RESET,WX6933);
	and 	XG17604 	(WX7167,RESET,WX6919);
	and 	XG17605 	(WX7165,RESET,WX6905);
	and 	XG17606 	(WX7163,RESET,WX6891);
	and 	XG17607 	(WX7161,RESET,WX6877);
	and 	XG17608 	(WX7159,RESET,WX6863);
	and 	XG17609 	(WX7157,RESET,WX6849);
	and 	XG17610 	(WX7155,RESET,WX6835);
	and 	XG17611 	(WX7153,RESET,WX6821);
	and 	XG17612 	(WX7151,RESET,WX6807);
	and 	XG17613 	(WX7149,RESET,WX6793);
	and 	XG17614 	(WX7147,RESET,WX6779);
	and 	XG17615 	(WX7145,RESET,WX6765);
	and 	XG17616 	(WX7143,RESET,WX6751);
	and 	XG17617 	(WX7141,RESET,WX6737);
	and 	XG17618 	(WX7139,RESET,WX6723);
	and 	XG17619 	(WX7137,RESET,WX6709);
	and 	XG17620 	(WX7135,RESET,WX6695);
	and 	XG17621 	(WX7133,RESET,WX6681);
	and 	XG17622 	(WX7131,RESET,WX6667);
	and 	XG17623 	(WX7129,RESET,WX6653);
	and 	XG17624 	(WX7127,RESET,WX6639);
	and 	XG17625 	(WX7125,RESET,WX6625);
	and 	XG17626 	(WX7123,RESET,WX6611);
	and 	XG17627 	(WX7121,RESET,WX6597);
	and 	XG17628 	(WX7119,RESET,WX6583);
	and 	XG17629 	(WX7117,RESET,WX6569);
	and 	XG17630 	(WX7115,RESET,WX6555);
	and 	XG17631 	(WX7113,RESET,WX6541);
	and 	XG17632 	(WX7111,RESET,WX6527);
	and 	XG17633 	(WX7109,RESET,WX6513);
	and 	XG17634 	(WX5878,RESET,WX5654);
	and 	XG17635 	(WX5876,RESET,WX5640);
	and 	XG17636 	(WX5874,RESET,WX5626);
	and 	XG17637 	(WX5872,RESET,WX5612);
	and 	XG17638 	(WX5870,RESET,WX5598);
	and 	XG17639 	(WX5868,RESET,WX5584);
	and 	XG17640 	(WX5866,RESET,WX5570);
	and 	XG17641 	(WX5864,RESET,WX5556);
	and 	XG17642 	(WX5862,RESET,WX5542);
	and 	XG17643 	(WX5860,RESET,WX5528);
	and 	XG17644 	(WX5858,RESET,WX5514);
	and 	XG17645 	(WX5856,RESET,WX5500);
	and 	XG17646 	(WX5854,RESET,WX5486);
	and 	XG17647 	(WX5852,RESET,WX5472);
	and 	XG17648 	(WX5850,RESET,WX5458);
	and 	XG17649 	(WX5848,RESET,WX5444);
	and 	XG17650 	(WX5846,RESET,WX5430);
	and 	XG17651 	(WX5844,RESET,WX5416);
	and 	XG17652 	(WX5842,RESET,WX5402);
	and 	XG17653 	(WX5840,RESET,WX5388);
	and 	XG17654 	(WX5838,RESET,WX5374);
	and 	XG17655 	(WX5836,RESET,WX5360);
	and 	XG17656 	(WX5834,RESET,WX5346);
	and 	XG17657 	(WX5832,RESET,WX5332);
	and 	XG17658 	(WX5830,RESET,WX5318);
	and 	XG17659 	(WX5828,RESET,WX5304);
	and 	XG17660 	(WX5826,RESET,WX5290);
	and 	XG17661 	(WX5824,RESET,WX5276);
	and 	XG17662 	(WX5822,RESET,WX5262);
	and 	XG17663 	(WX5820,RESET,WX5248);
	and 	XG17664 	(WX5818,RESET,WX5234);
	and 	XG17665 	(WX5816,RESET,WX5220);
	and 	XG17666 	(WX4585,RESET,WX4361);
	and 	XG17667 	(WX4583,RESET,WX4347);
	and 	XG17668 	(WX4581,RESET,WX4333);
	and 	XG17669 	(WX4579,RESET,WX4319);
	and 	XG17670 	(WX4577,RESET,WX4305);
	and 	XG17671 	(WX4575,RESET,WX4291);
	and 	XG17672 	(WX4573,RESET,WX4277);
	and 	XG17673 	(WX4571,RESET,WX4263);
	and 	XG17674 	(WX4569,RESET,WX4249);
	and 	XG17675 	(WX4567,RESET,WX4235);
	and 	XG17676 	(WX4565,RESET,WX4221);
	and 	XG17677 	(WX4563,RESET,WX4207);
	and 	XG17678 	(WX4561,RESET,WX4193);
	and 	XG17679 	(WX4559,RESET,WX4179);
	and 	XG17680 	(WX4557,RESET,WX4165);
	and 	XG17681 	(WX4555,RESET,WX4151);
	and 	XG17682 	(WX4553,RESET,WX4137);
	and 	XG17683 	(WX4551,RESET,WX4123);
	and 	XG17684 	(WX4549,RESET,WX4109);
	and 	XG17685 	(WX4547,RESET,WX4095);
	and 	XG17686 	(WX4545,RESET,WX4081);
	and 	XG17687 	(WX4543,RESET,WX4067);
	and 	XG17688 	(WX4541,RESET,WX4053);
	and 	XG17689 	(WX4539,RESET,WX4039);
	and 	XG17690 	(WX4537,RESET,WX4025);
	and 	XG17691 	(WX4535,RESET,WX4011);
	and 	XG17692 	(WX4533,RESET,WX3997);
	and 	XG17693 	(WX4531,RESET,WX3983);
	and 	XG17694 	(WX4529,RESET,WX3969);
	and 	XG17695 	(WX4527,RESET,WX3955);
	and 	XG17696 	(WX4525,RESET,WX3941);
	and 	XG17697 	(WX4523,RESET,WX3927);
	and 	XG17698 	(WX3292,RESET,WX3068);
	and 	XG17699 	(WX3290,RESET,WX3054);
	and 	XG17700 	(WX3288,RESET,WX3040);
	and 	XG17701 	(WX3286,RESET,WX3026);
	and 	XG17702 	(WX3284,RESET,WX3012);
	and 	XG17703 	(WX3282,RESET,WX2998);
	and 	XG17704 	(WX3280,RESET,WX2984);
	and 	XG17705 	(WX3278,RESET,WX2970);
	and 	XG17706 	(WX3276,RESET,WX2956);
	and 	XG17707 	(WX3274,RESET,WX2942);
	and 	XG17708 	(WX3272,RESET,WX2928);
	and 	XG17709 	(WX3270,RESET,WX2914);
	and 	XG17710 	(WX3268,RESET,WX2900);
	and 	XG17711 	(WX3266,RESET,WX2886);
	and 	XG17712 	(WX3264,RESET,WX2872);
	and 	XG17713 	(WX3262,RESET,WX2858);
	and 	XG17714 	(WX3260,RESET,WX2844);
	and 	XG17715 	(WX3258,RESET,WX2830);
	and 	XG17716 	(WX3256,RESET,WX2816);
	and 	XG17717 	(WX3254,RESET,WX2802);
	and 	XG17718 	(WX3252,RESET,WX2788);
	and 	XG17719 	(WX3250,RESET,WX2774);
	and 	XG17720 	(WX3248,RESET,WX2760);
	and 	XG17721 	(WX3246,RESET,WX2746);
	and 	XG17722 	(WX3244,RESET,WX2732);
	and 	XG17723 	(WX3242,RESET,WX2718);
	and 	XG17724 	(WX3240,RESET,WX2704);
	and 	XG17725 	(WX3238,RESET,WX2690);
	and 	XG17726 	(WX3236,RESET,WX2676);
	and 	XG17727 	(WX3234,RESET,WX2662);
	and 	XG17728 	(WX3232,RESET,WX2648);
	and 	XG17729 	(WX3230,RESET,WX2634);
	and 	XG17730 	(WX1999,RESET,WX1775);
	and 	XG17731 	(WX1997,RESET,WX1761);
	and 	XG17732 	(WX1995,RESET,WX1747);
	and 	XG17733 	(WX1993,RESET,WX1733);
	and 	XG17734 	(WX1991,RESET,WX1719);
	and 	XG17735 	(WX1989,RESET,WX1705);
	and 	XG17736 	(WX1987,RESET,WX1691);
	and 	XG17737 	(WX1985,RESET,WX1677);
	and 	XG17738 	(WX1983,RESET,WX1663);
	and 	XG17739 	(WX1981,RESET,WX1649);
	and 	XG17740 	(WX1979,RESET,WX1635);
	and 	XG17741 	(WX1977,RESET,WX1621);
	and 	XG17742 	(WX1975,RESET,WX1607);
	and 	XG17743 	(WX1973,RESET,WX1593);
	and 	XG17744 	(WX1971,RESET,WX1579);
	and 	XG17745 	(WX1969,RESET,WX1565);
	and 	XG17746 	(WX1967,RESET,WX1551);
	and 	XG17747 	(WX1965,RESET,WX1537);
	and 	XG17748 	(WX1963,RESET,WX1523);
	and 	XG17749 	(WX1961,RESET,WX1509);
	and 	XG17750 	(WX1959,RESET,WX1495);
	and 	XG17751 	(WX1957,RESET,WX1481);
	and 	XG17752 	(WX1955,RESET,WX1467);
	and 	XG17753 	(WX1953,RESET,WX1453);
	and 	XG17754 	(WX1951,RESET,WX1439);
	and 	XG17755 	(WX1949,RESET,WX1425);
	and 	XG17756 	(WX1947,RESET,WX1411);
	and 	XG17757 	(WX1945,RESET,WX1397);
	and 	XG17758 	(WX1943,RESET,WX1383);
	and 	XG17759 	(WX1941,RESET,WX1369);
	and 	XG17760 	(WX1939,RESET,WX1355);
	and 	XG17761 	(WX1937,RESET,WX1341);
	and 	XG17762 	(WX706,RESET,WX482);
	and 	XG17763 	(WX704,RESET,WX468);
	and 	XG17764 	(WX702,RESET,WX454);
	and 	XG17765 	(WX700,RESET,WX440);
	and 	XG17766 	(WX698,RESET,WX426);
	and 	XG17767 	(WX696,RESET,WX412);
	and 	XG17768 	(WX694,RESET,WX398);
	and 	XG17769 	(WX692,RESET,WX384);
	and 	XG17770 	(WX690,RESET,WX370);
	and 	XG17771 	(WX688,RESET,WX356);
	and 	XG17772 	(WX686,RESET,WX342);
	and 	XG17773 	(WX684,RESET,WX328);
	and 	XG17774 	(WX682,RESET,WX314);
	and 	XG17775 	(WX680,RESET,WX300);
	and 	XG17776 	(WX678,RESET,WX286);
	and 	XG17777 	(WX676,RESET,WX272);
	and 	XG17778 	(WX674,RESET,WX258);
	and 	XG17779 	(WX672,RESET,WX244);
	and 	XG17780 	(WX670,RESET,WX230);
	and 	XG17781 	(WX668,RESET,WX216);
	and 	XG17782 	(WX666,RESET,WX202);
	and 	XG17783 	(WX664,RESET,WX188);
	and 	XG17784 	(WX662,RESET,WX174);
	and 	XG17785 	(WX660,RESET,WX160);
	and 	XG17786 	(WX658,RESET,WX146);
	and 	XG17787 	(WX656,RESET,WX132);
	and 	XG17788 	(WX654,RESET,WX118);
	and 	XG17789 	(WX652,RESET,WX104);
	and 	XG17790 	(WX650,RESET,WX90);
	and 	XG17791 	(WX648,RESET,WX76);
	and 	XG17792 	(WX646,RESET,WX62);
	and 	XG17793 	(WX644,RESET,WX48);
	not 	XG17794 	(DATA_9_31,WX1011);
	not 	XG17795 	(DATA_9_30,WX1018);
	not 	XG17796 	(DATA_9_29,WX1025);
	not 	XG17797 	(DATA_9_28,WX1032);
	not 	XG17798 	(DATA_9_27,WX1039);
	not 	XG17799 	(DATA_9_26,WX1046);
	not 	XG17800 	(DATA_9_25,WX1053);
	not 	XG17801 	(DATA_9_24,WX1060);
	not 	XG17802 	(DATA_9_23,WX1067);
	not 	XG17803 	(DATA_9_22,WX1074);
	not 	XG17804 	(DATA_9_21,WX1081);
	not 	XG17805 	(DATA_9_20,WX1088);
	not 	XG17806 	(DATA_9_19,WX1095);
	not 	XG17807 	(DATA_9_18,WX1102);
	not 	XG17808 	(DATA_9_17,WX1109);
	not 	XG17809 	(DATA_9_16,WX1116);
	not 	XG17810 	(DATA_9_15,WX1123);
	not 	XG17811 	(DATA_9_14,WX1130);
	not 	XG17812 	(DATA_9_13,WX1137);
	not 	XG17813 	(DATA_9_12,WX1144);
	not 	XG17814 	(DATA_9_11,WX1151);
	not 	XG17815 	(DATA_9_10,WX1158);
	not 	XG17816 	(DATA_9_9,WX1165);
	not 	XG17817 	(DATA_9_8,WX1172);
	not 	XG17818 	(DATA_9_7,WX1179);
	not 	XG17819 	(DATA_9_6,WX1186);
	not 	XG17820 	(DATA_9_5,WX1193);
	not 	XG17821 	(DATA_9_4,WX1200);
	not 	XG17822 	(DATA_9_3,WX1207);
	not 	XG17823 	(DATA_9_2,WX1214);
	not 	XG17824 	(DATA_9_1,WX1221);
	not 	XG17825 	(DATA_9_0,WX1228);
	dff 	XG17826 	(CRC_OUT_9_0,WX1264);
	dff 	XG17827 	(CRC_OUT_9_1,WX1266);
	dff 	XG17828 	(CRC_OUT_9_2,WX1268);
	dff 	XG17829 	(CRC_OUT_9_3,WX1270);
	dff 	XG17830 	(CRC_OUT_9_4,WX1272);
	dff 	XG17831 	(CRC_OUT_9_5,WX1274);
	dff 	XG17832 	(CRC_OUT_9_6,WX1276);
	dff 	XG17833 	(CRC_OUT_9_7,WX1278);
	dff 	XG17834 	(CRC_OUT_9_8,WX1280);
	dff 	XG17835 	(CRC_OUT_9_9,WX1282);
	dff 	XG17836 	(CRC_OUT_9_10,WX1284);
	dff 	XG17837 	(CRC_OUT_9_11,WX1286);
	dff 	XG17838 	(CRC_OUT_9_12,WX1288);
	dff 	XG17839 	(CRC_OUT_9_13,WX1290);
	dff 	XG17840 	(CRC_OUT_9_14,WX1292);
	dff 	XG17841 	(CRC_OUT_9_15,WX1294);
	dff 	XG17842 	(CRC_OUT_9_16,WX1296);
	dff 	XG17843 	(CRC_OUT_9_17,WX1298);
	dff 	XG17844 	(CRC_OUT_9_18,WX1300);
	dff 	XG17845 	(CRC_OUT_9_19,WX1302);
	dff 	XG17846 	(CRC_OUT_9_20,WX1304);
	dff 	XG17847 	(CRC_OUT_9_21,WX1306);
	dff 	XG17848 	(CRC_OUT_9_22,WX1308);
	dff 	XG17849 	(CRC_OUT_9_23,WX1310);
	dff 	XG17850 	(CRC_OUT_9_24,WX1312);
	dff 	XG17851 	(CRC_OUT_9_25,WX1314);
	dff 	XG17852 	(CRC_OUT_9_26,WX1316);
	dff 	XG17853 	(CRC_OUT_9_27,WX1318);
	dff 	XG17854 	(CRC_OUT_9_28,WX1320);
	dff 	XG17855 	(CRC_OUT_9_29,WX1322);
	dff 	XG17856 	(CRC_OUT_9_30,WX1324);
	dff 	XG17857 	(CRC_OUT_9_31,WX1326);
	dff 	XG17858 	(CRC_OUT_8_0,WX2557);
	dff 	XG17859 	(CRC_OUT_8_1,WX2559);
	dff 	XG17860 	(CRC_OUT_8_2,WX2561);
	dff 	XG17861 	(CRC_OUT_8_3,WX2563);
	dff 	XG17862 	(CRC_OUT_8_4,WX2565);
	dff 	XG17863 	(CRC_OUT_8_5,WX2567);
	dff 	XG17864 	(CRC_OUT_8_6,WX2569);
	dff 	XG17865 	(CRC_OUT_8_7,WX2571);
	dff 	XG17866 	(CRC_OUT_8_8,WX2573);
	dff 	XG17867 	(CRC_OUT_8_9,WX2575);
	dff 	XG17868 	(CRC_OUT_8_10,WX2577);
	dff 	XG17869 	(CRC_OUT_8_11,WX2579);
	dff 	XG17870 	(CRC_OUT_8_12,WX2581);
	dff 	XG17871 	(CRC_OUT_8_13,WX2583);
	dff 	XG17872 	(CRC_OUT_8_14,WX2585);
	dff 	XG17873 	(CRC_OUT_8_15,WX2587);
	dff 	XG17874 	(CRC_OUT_8_16,WX2589);
	dff 	XG17875 	(CRC_OUT_8_17,WX2591);
	dff 	XG17876 	(CRC_OUT_8_18,WX2593);
	dff 	XG17877 	(CRC_OUT_8_19,WX2595);
	dff 	XG17878 	(CRC_OUT_8_20,WX2597);
	dff 	XG17879 	(CRC_OUT_8_21,WX2599);
	dff 	XG17880 	(CRC_OUT_8_22,WX2601);
	dff 	XG17881 	(CRC_OUT_8_23,WX2603);
	dff 	XG17882 	(CRC_OUT_8_24,WX2605);
	dff 	XG17883 	(CRC_OUT_8_25,WX2607);
	dff 	XG17884 	(CRC_OUT_8_26,WX2609);
	dff 	XG17885 	(CRC_OUT_8_27,WX2611);
	dff 	XG17886 	(CRC_OUT_8_28,WX2613);
	dff 	XG17887 	(CRC_OUT_8_29,WX2615);
	dff 	XG17888 	(CRC_OUT_8_30,WX2617);
	dff 	XG17889 	(CRC_OUT_8_31,WX2619);
	dff 	XG17890 	(CRC_OUT_7_0,WX3850);
	dff 	XG17891 	(CRC_OUT_7_1,WX3852);
	dff 	XG17892 	(CRC_OUT_7_2,WX3854);
	dff 	XG17893 	(CRC_OUT_7_3,WX3856);
	dff 	XG17894 	(CRC_OUT_7_4,WX3858);
	dff 	XG17895 	(CRC_OUT_7_5,WX3860);
	dff 	XG17896 	(CRC_OUT_7_6,WX3862);
	dff 	XG17897 	(CRC_OUT_7_7,WX3864);
	dff 	XG17898 	(CRC_OUT_7_8,WX3866);
	dff 	XG17899 	(CRC_OUT_7_9,WX3868);
	dff 	XG17900 	(CRC_OUT_7_10,WX3870);
	dff 	XG17901 	(CRC_OUT_7_11,WX3872);
	dff 	XG17902 	(CRC_OUT_7_12,WX3874);
	dff 	XG17903 	(CRC_OUT_7_13,WX3876);
	dff 	XG17904 	(CRC_OUT_7_14,WX3878);
	dff 	XG17905 	(CRC_OUT_7_15,WX3880);
	dff 	XG17906 	(CRC_OUT_7_16,WX3882);
	dff 	XG17907 	(CRC_OUT_7_17,WX3884);
	dff 	XG17908 	(CRC_OUT_7_18,WX3886);
	dff 	XG17909 	(CRC_OUT_7_19,WX3888);
	dff 	XG17910 	(CRC_OUT_7_20,WX3890);
	dff 	XG17911 	(CRC_OUT_7_21,WX3892);
	dff 	XG17912 	(CRC_OUT_7_22,WX3894);
	dff 	XG17913 	(CRC_OUT_7_23,WX3896);
	dff 	XG17914 	(CRC_OUT_7_24,WX3898);
	dff 	XG17915 	(CRC_OUT_7_25,WX3900);
	dff 	XG17916 	(CRC_OUT_7_26,WX3902);
	dff 	XG17917 	(CRC_OUT_7_27,WX3904);
	dff 	XG17918 	(CRC_OUT_7_28,WX3906);
	dff 	XG17919 	(CRC_OUT_7_29,WX3908);
	dff 	XG17920 	(CRC_OUT_7_30,WX3910);
	dff 	XG17921 	(CRC_OUT_7_31,WX3912);
	dff 	XG17922 	(CRC_OUT_6_0,WX5143);
	dff 	XG17923 	(CRC_OUT_6_1,WX5145);
	dff 	XG17924 	(CRC_OUT_6_2,WX5147);
	dff 	XG17925 	(CRC_OUT_6_3,WX5149);
	dff 	XG17926 	(CRC_OUT_6_4,WX5151);
	dff 	XG17927 	(CRC_OUT_6_5,WX5153);
	dff 	XG17928 	(CRC_OUT_6_6,WX5155);
	dff 	XG17929 	(CRC_OUT_6_7,WX5157);
	dff 	XG17930 	(CRC_OUT_6_8,WX5159);
	dff 	XG17931 	(CRC_OUT_6_9,WX5161);
	dff 	XG17932 	(CRC_OUT_6_10,WX5163);
	dff 	XG17933 	(CRC_OUT_6_11,WX5165);
	dff 	XG17934 	(CRC_OUT_6_12,WX5167);
	dff 	XG17935 	(CRC_OUT_6_13,WX5169);
	dff 	XG17936 	(CRC_OUT_6_14,WX5171);
	dff 	XG17937 	(CRC_OUT_6_15,WX5173);
	dff 	XG17938 	(CRC_OUT_6_16,WX5175);
	dff 	XG17939 	(CRC_OUT_6_17,WX5177);
	dff 	XG17940 	(CRC_OUT_6_18,WX5179);
	dff 	XG17941 	(CRC_OUT_6_19,WX5181);
	dff 	XG17942 	(CRC_OUT_6_20,WX5183);
	dff 	XG17943 	(CRC_OUT_6_21,WX5185);
	dff 	XG17944 	(CRC_OUT_6_22,WX5187);
	dff 	XG17945 	(CRC_OUT_6_23,WX5189);
	dff 	XG17946 	(CRC_OUT_6_24,WX5191);
	dff 	XG17947 	(CRC_OUT_6_25,WX5193);
	dff 	XG17948 	(CRC_OUT_6_26,WX5195);
	dff 	XG17949 	(CRC_OUT_6_27,WX5197);
	dff 	XG17950 	(CRC_OUT_6_28,WX5199);
	dff 	XG17951 	(CRC_OUT_6_29,WX5201);
	dff 	XG17952 	(CRC_OUT_6_30,WX5203);
	dff 	XG17953 	(CRC_OUT_6_31,WX5205);
	dff 	XG17954 	(CRC_OUT_5_0,WX6436);
	dff 	XG17955 	(CRC_OUT_5_1,WX6438);
	dff 	XG17956 	(CRC_OUT_5_2,WX6440);
	dff 	XG17957 	(CRC_OUT_5_3,WX6442);
	dff 	XG17958 	(CRC_OUT_5_4,WX6444);
	dff 	XG17959 	(CRC_OUT_5_5,WX6446);
	dff 	XG17960 	(CRC_OUT_5_6,WX6448);
	dff 	XG17961 	(CRC_OUT_5_7,WX6450);
	dff 	XG17962 	(CRC_OUT_5_8,WX6452);
	dff 	XG17963 	(CRC_OUT_5_9,WX6454);
	dff 	XG17964 	(CRC_OUT_5_10,WX6456);
	dff 	XG17965 	(CRC_OUT_5_11,WX6458);
	dff 	XG17966 	(CRC_OUT_5_12,WX6460);
	dff 	XG17967 	(CRC_OUT_5_13,WX6462);
	dff 	XG17968 	(CRC_OUT_5_14,WX6464);
	dff 	XG17969 	(CRC_OUT_5_15,WX6466);
	dff 	XG17970 	(CRC_OUT_5_16,WX6468);
	dff 	XG17971 	(CRC_OUT_5_17,WX6470);
	dff 	XG17972 	(CRC_OUT_5_18,WX6472);
	dff 	XG17973 	(CRC_OUT_5_19,WX6474);
	dff 	XG17974 	(CRC_OUT_5_20,WX6476);
	dff 	XG17975 	(CRC_OUT_5_21,WX6478);
	dff 	XG17976 	(CRC_OUT_5_22,WX6480);
	dff 	XG17977 	(CRC_OUT_5_23,WX6482);
	dff 	XG17978 	(CRC_OUT_5_24,WX6484);
	dff 	XG17979 	(CRC_OUT_5_25,WX6486);
	dff 	XG17980 	(CRC_OUT_5_26,WX6488);
	dff 	XG17981 	(CRC_OUT_5_27,WX6490);
	dff 	XG17982 	(CRC_OUT_5_28,WX6492);
	dff 	XG17983 	(CRC_OUT_5_29,WX6494);
	dff 	XG17984 	(CRC_OUT_5_30,WX6496);
	dff 	XG17985 	(CRC_OUT_5_31,WX6498);
	dff 	XG17986 	(CRC_OUT_4_0,WX7729);
	dff 	XG17987 	(CRC_OUT_4_1,WX7731);
	dff 	XG17988 	(CRC_OUT_4_2,WX7733);
	dff 	XG17989 	(CRC_OUT_4_3,WX7735);
	dff 	XG17990 	(CRC_OUT_4_4,WX7737);
	dff 	XG17991 	(CRC_OUT_4_5,WX7739);
	dff 	XG17992 	(CRC_OUT_4_6,WX7741);
	dff 	XG17993 	(CRC_OUT_4_7,WX7743);
	dff 	XG17994 	(CRC_OUT_4_8,WX7745);
	dff 	XG17995 	(CRC_OUT_4_9,WX7747);
	dff 	XG17996 	(CRC_OUT_4_10,WX7749);
	dff 	XG17997 	(CRC_OUT_4_11,WX7751);
	dff 	XG17998 	(CRC_OUT_4_12,WX7753);
	dff 	XG17999 	(CRC_OUT_4_13,WX7755);
	dff 	XG18000 	(CRC_OUT_4_14,WX7757);
	dff 	XG18001 	(CRC_OUT_4_15,WX7759);
	dff 	XG18002 	(CRC_OUT_4_16,WX7761);
	dff 	XG18003 	(CRC_OUT_4_17,WX7763);
	dff 	XG18004 	(CRC_OUT_4_18,WX7765);
	dff 	XG18005 	(CRC_OUT_4_19,WX7767);
	dff 	XG18006 	(CRC_OUT_4_20,WX7769);
	dff 	XG18007 	(CRC_OUT_4_21,WX7771);
	dff 	XG18008 	(CRC_OUT_4_22,WX7773);
	dff 	XG18009 	(CRC_OUT_4_23,WX7775);
	dff 	XG18010 	(CRC_OUT_4_24,WX7777);
	dff 	XG18011 	(CRC_OUT_4_25,WX7779);
	dff 	XG18012 	(CRC_OUT_4_26,WX7781);
	dff 	XG18013 	(CRC_OUT_4_27,WX7783);
	dff 	XG18014 	(CRC_OUT_4_28,WX7785);
	dff 	XG18015 	(CRC_OUT_4_29,WX7787);
	dff 	XG18016 	(CRC_OUT_4_30,WX7789);
	dff 	XG18017 	(CRC_OUT_4_31,WX7791);
	dff 	XG18018 	(CRC_OUT_3_0,WX9022);
	dff 	XG18019 	(CRC_OUT_3_1,WX9024);
	dff 	XG18020 	(CRC_OUT_3_2,WX9026);
	dff 	XG18021 	(CRC_OUT_3_3,WX9028);
	dff 	XG18022 	(CRC_OUT_3_4,WX9030);
	dff 	XG18023 	(CRC_OUT_3_5,WX9032);
	dff 	XG18024 	(CRC_OUT_3_6,WX9034);
	dff 	XG18025 	(CRC_OUT_3_7,WX9036);
	dff 	XG18026 	(CRC_OUT_3_8,WX9038);
	dff 	XG18027 	(CRC_OUT_3_9,WX9040);
	dff 	XG18028 	(CRC_OUT_3_10,WX9042);
	dff 	XG18029 	(CRC_OUT_3_11,WX9044);
	dff 	XG18030 	(CRC_OUT_3_12,WX9046);
	dff 	XG18031 	(CRC_OUT_3_13,WX9048);
	dff 	XG18032 	(CRC_OUT_3_14,WX9050);
	dff 	XG18033 	(CRC_OUT_3_15,WX9052);
	dff 	XG18034 	(CRC_OUT_3_16,WX9054);
	dff 	XG18035 	(CRC_OUT_3_17,WX9056);
	dff 	XG18036 	(CRC_OUT_3_18,WX9058);
	dff 	XG18037 	(CRC_OUT_3_19,WX9060);
	dff 	XG18038 	(CRC_OUT_3_20,WX9062);
	dff 	XG18039 	(CRC_OUT_3_21,WX9064);
	dff 	XG18040 	(CRC_OUT_3_22,WX9066);
	dff 	XG18041 	(CRC_OUT_3_23,WX9068);
	dff 	XG18042 	(CRC_OUT_3_24,WX9070);
	dff 	XG18043 	(CRC_OUT_3_25,WX9072);
	dff 	XG18044 	(CRC_OUT_3_26,WX9074);
	dff 	XG18045 	(CRC_OUT_3_27,WX9076);
	dff 	XG18046 	(CRC_OUT_3_28,WX9078);
	dff 	XG18047 	(CRC_OUT_3_29,WX9080);
	dff 	XG18048 	(CRC_OUT_3_30,WX9082);
	dff 	XG18049 	(CRC_OUT_3_31,WX9084);
	dff 	XG18050 	(CRC_OUT_2_0,WX10315);
	dff 	XG18051 	(CRC_OUT_2_1,WX10317);
	dff 	XG18052 	(CRC_OUT_2_2,WX10319);
	dff 	XG18053 	(CRC_OUT_2_3,WX10321);
	dff 	XG18054 	(CRC_OUT_2_4,WX10323);
	dff 	XG18055 	(CRC_OUT_2_5,WX10325);
	dff 	XG18056 	(CRC_OUT_2_6,WX10327);
	dff 	XG18057 	(CRC_OUT_2_7,WX10329);
	dff 	XG18058 	(CRC_OUT_2_8,WX10331);
	dff 	XG18059 	(CRC_OUT_2_9,WX10333);
	dff 	XG18060 	(CRC_OUT_2_10,WX10335);
	dff 	XG18061 	(CRC_OUT_2_11,WX10337);
	dff 	XG18062 	(CRC_OUT_2_12,WX10339);
	dff 	XG18063 	(CRC_OUT_2_13,WX10341);
	dff 	XG18064 	(CRC_OUT_2_14,WX10343);
	dff 	XG18065 	(CRC_OUT_2_15,WX10345);
	dff 	XG18066 	(CRC_OUT_2_16,WX10347);
	dff 	XG18067 	(CRC_OUT_2_17,WX10349);
	dff 	XG18068 	(CRC_OUT_2_18,WX10351);
	dff 	XG18069 	(CRC_OUT_2_19,WX10353);
	dff 	XG18070 	(CRC_OUT_2_20,WX10355);
	dff 	XG18071 	(CRC_OUT_2_21,WX10357);
	dff 	XG18072 	(CRC_OUT_2_22,WX10359);
	dff 	XG18073 	(CRC_OUT_2_23,WX10361);
	dff 	XG18074 	(CRC_OUT_2_24,WX10363);
	dff 	XG18075 	(CRC_OUT_2_25,WX10365);
	dff 	XG18076 	(CRC_OUT_2_26,WX10367);
	dff 	XG18077 	(CRC_OUT_2_27,WX10369);
	dff 	XG18078 	(CRC_OUT_2_28,WX10371);
	dff 	XG18079 	(CRC_OUT_2_29,WX10373);
	dff 	XG18080 	(CRC_OUT_2_30,WX10375);
	dff 	XG18081 	(CRC_OUT_2_31,WX10377);
	dff 	XG18082 	(CRC_OUT_1_0,WX11608);
	dff 	XG18083 	(CRC_OUT_1_1,WX11610);
	dff 	XG18084 	(CRC_OUT_1_2,WX11612);
	dff 	XG18085 	(CRC_OUT_1_3,WX11614);
	dff 	XG18086 	(CRC_OUT_1_4,WX11616);
	dff 	XG18087 	(CRC_OUT_1_5,WX11618);
	dff 	XG18088 	(CRC_OUT_1_6,WX11620);
	dff 	XG18089 	(CRC_OUT_1_7,WX11622);
	dff 	XG18090 	(CRC_OUT_1_8,WX11624);
	dff 	XG18091 	(CRC_OUT_1_9,WX11626);
	dff 	XG18092 	(CRC_OUT_1_10,WX11628);
	dff 	XG18093 	(CRC_OUT_1_11,WX11630);
	dff 	XG18094 	(CRC_OUT_1_12,WX11632);
	dff 	XG18095 	(CRC_OUT_1_13,WX11634);
	dff 	XG18096 	(CRC_OUT_1_14,WX11636);
	dff 	XG18097 	(CRC_OUT_1_15,WX11638);
	dff 	XG18098 	(CRC_OUT_1_16,WX11640);
	dff 	XG18099 	(CRC_OUT_1_17,WX11642);
	dff 	XG18100 	(CRC_OUT_1_18,WX11644);
	dff 	XG18101 	(CRC_OUT_1_19,WX11646);
	dff 	XG18102 	(CRC_OUT_1_20,WX11648);
	dff 	XG18103 	(CRC_OUT_1_21,WX11650);
	dff 	XG18104 	(CRC_OUT_1_22,WX11652);
	dff 	XG18105 	(CRC_OUT_1_23,WX11654);
	dff 	XG18106 	(CRC_OUT_1_24,WX11656);
	dff 	XG18107 	(CRC_OUT_1_25,WX11658);
	dff 	XG18108 	(CRC_OUT_1_26,WX11660);
	dff 	XG18109 	(CRC_OUT_1_27,WX11662);
	dff 	XG18110 	(CRC_OUT_1_28,WX11664);
	dff 	XG18111 	(CRC_OUT_1_29,WX11666);
	dff 	XG18112 	(CRC_OUT_1_30,WX11668);
	dff 	XG18113 	(CRC_OUT_1_31,WX11670);

endmodule
