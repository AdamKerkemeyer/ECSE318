--VHDL
