--Traffic Light Controller